-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǑ[�������n� �2��2�������T��_�[���n� �0���s�"���0����wH��[Uװ���!�u�g��n�d����������h��A��
�u�&�2�9�/����Y����wF�N��U���u�<�!�2�%�g�W��Y����f+��c/��U���u�<�!�2�%�g�W��Y����Z��`'��=���u�u�o�;�2�8�W��J��ƹF��^ ��"����u�u�u�m�3����Y���]ǻN��������u�w�}�M�������	[�UךU���<�a����}�W���C����T��S��G�ߊu�u�<�`� ��?���Y���Z��P��O���g�_�u�u�>�k� ���1���F�^ �����o�u�g�_�w�}����.����F�N�����2�'�o�u�e�W�W����ޓ�z"��N��U���<�!�2�'�m�}�E�ԜY�ƨ�]_��~*��U���u�u�<�!�0�/�M���K���F��Y_��"����u�u�u�m�3����Y���]ǻN����
���u�w�}�Wշ�����\�\�U���1�;�g����W���Y�ܥ�G��EN�U��_�u�u�<�f��>���Y���F��Y�����h�f�n�u�w�9����.����F�N�����2�'�o�u�e�W�W�������d/��N��U���o�;�0�0�w�`�D��Y����Z��h9��!���u�u�u�<�#�:���Y����F�S��B�����u�u�w�g��������U��=N��U���!����w�}�W�������V�
N�\���:�!�}�u�w�9����Yɏ����h�����0�!�'�d�w�2����I��ƹF��^ �U���;�u�!�
�8�4�(������F��@ ��U���_�u�u�<�d�}�M���Y����_	��T1�����}�`�1�"�#�}�^�ԜY�ƨ�]R�T��Uʦ�1�9�2�6�!�>����Lӂ��]��G�U���1�;�u�u�>�}��������l��C��D���:�;�:�e�l�}�WϺ����	����*���<�
�0�!�%�l�W������]ǻN����u�o�;�u�#�����&����\�N�����u�|�_�u�w�4�O���C���@��[�����6�:�}�`�3�*����P���F��YW��Uм�u�&�1�9�0�>����������Y��E��u�u�1�;�g�}�M���Y����_	��T1�����}�`�1�"�#�}�^�ԜY�ƨ�]W��N�����!�
�:�<��8����H�ƨ�D��^����u�<�d�u�w�4�Wϭ�����Z��R����u�:�;�:�g�f�W�������F�^ �����9�2�6�#�4�2�_������\F��d��Uʱ�;�a�u�o�9�}��������E��X��@ʱ�"�!�u�|�]�}�W���H���	����*���<�
�0�!�%�l�W������]ǻN����u�u�<�u�$�9��������G	��[�����:�e�n�u�w�9���Y�ܥ�F��S1�����#�6�:�}�w�2����I��ƹF��X��U���o� �u�!��2��������W��S�����|�n�0�1�2�)���s����Z��C��U���u�3�8��f��3���&����P��1��ފ�c�d�<�_�w�}�ZϮ��ƥ�G��V�����9�_�u�u�>�3�ϭ����	F��S1�����#�6�:�}�w�2����I��ƹF�N�����d�&�2�4�$�}�Wϭ�����^��1�U���u�!�
�:�>���������W	��C��\�ߊu�u�<�;�;�0����H���	F��S1�����#�6�:�}�b�9� ���Y����F�D����� �
�
�u�w�g��������l��C��D���:�;�:�e�l�}�Wϭ�����^��1�U���u�!�
�:�>���������W	��C��\�ߊu�u�<�;�;�0����M���	F��S1�����#�6�:�}�b�9� ���Y����F�D����� �
�
�u�w�g��������l��C��D���:�;�:�e�l�}�Wϭ�����^��1�U���u�!�
�:�>���������W	��C��\�ߊu�u�<�;�;�0����N���	F��S1�����#�6�:�}�b�9� ���Y����F�C�����u�u�<�;�;�W�W���������h\��U���o�&�1�9�0�>����������Y��E��u�u�&�2�6�}����&���\��C
�����
�0�!�'�f�}�������9F������8�-�g�g�w�}�W���&����P9��T��]���1�"�!�u�~�W�W���������h\��U���o�&�1�9�0�>����������Y��E��u�u�x�u�2�8�W�������@l�N�����u� �
�
�w�}�Mϭ�����Z��R����u�:�;�:�g�f�W���
����_F��O1��D���u�u�!�
�8�4�(������F��@ ��U���_�u�u�x�;�+���
����_ǻN�����9�8�-�a�g�}�W�������T��A�����`�1�"�!�w�t�}�������V
�
N����_�x�u�0�2�<�ϲ����
��^�� ���
�u�h�1�9�}����
���F�^�����u�<�g�_�"��(���Dӂ�� F��R �����|�h�r�r�2�.�W���M���K9��N�U���`�"�0�u�2�u�^��^����_��S��N��-�d�f�i�w�4�@ϩ��ƿ�_N��S��E���9�0�1�;�l�0����M���W����ʦ�9�e�u�u�g�}��������l��O1��@��u�<�d�u�?�3����I���V�R��U���d�n�8�-�f�k�K�������D����]���h�r�r�0�$�}���B����lW��R�����`�"�0�u�2�u�^��^����_��S��C�ߠx�u�0�0�6�8��������\��=��*؊�u�h�8�-�f�m� ���Y����O�I�U���0�8�-�d�f�W����&�����h_��U���;�&�9�d�w�}�G�������F��h]����g�g�i�u�"��(�������V
�N��R��0�&�u� ���L���ԓ�Z�Z��D��"�0�u�0��t�J���^Ӄ��VF��O1��B�ߠx�u�0�0�6�8��������\��=��*ي�u�h�8�-�e�m� ���Y����O�I�U���0�8�-�g�f�W����&�����h\��U���;�&�9�g�w�}�G�������F��h]�����;�'�!�w�8����Y����Pl��O1��E��u� �
�
�w�5�ϭ����F�N����� �
�
�n�]�p�����Ơ�T��S��U��8�-�a�e�]�8�Ͽ�����P��RU�