-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��l����}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���_�u�u�
����������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��V�����u������4�ԜY�Ƽ�9��N��U���
���
��	�%���Lӂ��]��G�U���%�e�g�4��1�W���7ӵ��l*��~-�U���%�e�f�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I�Փ�C9��SN�<����
���l�}�WϮ�I���/��d:��9�������w�l�W������]ǻN��*ڊ�
�%�#�1�m��W���&����p]ǻN��*ڊ�u�u�����0���/����aF�N�����u�|�_�u�w��(ځ�	����\��yN��1�����_�u�w��(���Y����g"��x)��*�����}�`�3�*����P���F��1�����9�u�u����;���:���F��1�Oʜ�u��
����2���+������Y��E��u�u�%�e�`�<�(���Y�ƅ�5��h"��<��u�u�%�e�o�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӖ��l^��G1�����u��
���L���YӖ��l_�'��&���������W��Y����G	�UךU���
�
�
�%�!�9�Mϗ�Y����)��tUךU���
�
�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I����R��[
��U��������W�W���&ù��\��yN��1��������}�F�������V�=N��U���
�d�4�
�;�}�W���*����|!��d��Uʥ�e�d�u�u���3���>����v%��eN��@ʱ�"�!�u�|�]�}�W���&�ԓ�C9��SN�<����
���l�}�WϮ�I����	F��=��*����
����u�BϺ�����O��N�����d�
�%�#�3�g�>���-����t/��=N��U���
�a�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����Hǹ��l��T��;ʆ�����]�}�W���&���/��d:��9�������w�l�W������]ǻN��*ڊ�`�4�
�9�w�}�9ύ�=����z%��N����o��u����>���<����N��
�����e�n�u�u�'�l��������z(��c*��:���n�u�u�%�b�m�Mϗ�Y����)��t1��6���u�d�u�:�9�2�G��Y����lS��h�����o��u����>��Y����lS��T��;ʆ�������8���H�ƨ�D��^����u�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�u�w��$���5����l0��c!��]���1�"�!�u�~�W�W���&ƹ��R��[
��U��������W�W���&ƹ��	F��=��*����
����u�BϺ�����O��N�����f�4�
�9�w�}�9ύ�=����z%��N�����a�o��u���8���&����|4�[�����:�e�n�u�w�-�B�������WF��~ ��!�����n�u�w�-�B��Cӯ��`2��{!��6�����u�d�w�2����I��ƹF��h[��*���#�1�o��w�	�(���0��ƹF��h[��U���������!���6���F��@ ��U���_�u�u�
����������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��V�����u������4�ԜY�Ƽ�9��N��U���
���
��	�%���Lӂ��]��G�U���%�`�m�4��1�W���7ӵ��l*��~-�U���%�`�l�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�L�ߓ�C9��SN�<����
���l�}�WϮ�L����	F��=��*����
����u�BϺ�����O��N�����d�
�%�#�3�g�>���-����t/��=N��U���
�d�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����H¹��l��T��;ʆ�����]�}�W���&���/��d:��9�������w�l�W������]ǻN��*ߊ�g�4�
�9�w�}�9ύ�=����z%��N�����d�u�u����;���:����g)��_����!�u�|�_�w�}�(ځ�J����E
��N��U���
���n�w�}����H����z(��c*��:���
�����h��������l�N��@��
�%�#�1�m��W���&����p]ǻN��*ߊ�`�o��u���8���&����|4�[�����:�e�n�u�w�-�B��&����_�'��&������_�w�}�(؁�Y�ƅ�5��h"��<������}�b�9� ���Y����F�G1��E���
�9�u�u���3���>����F�G1��D���u��
���(���-���S��X����n�u�u�%�`�l��������z(��c*��:���n�u�u�%�`�o�Mϗ�Y����)��t1��6���u�d�u�:�9�2�G��Y����lQ��h�����o��u����>��Y����lQ��T��;ʆ�������8���H�ƨ�D��^����u�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�u�w��$���5����l0��c!��]���1�"�!�u�~�W�W���&Ĺ��R��[
��U��������W�W���&Ĺ��	F��=��*����
����u�BϺ�����O��N�����`�4�
�9�w�}�9ύ�=����z%��N�����c�o��u���8���&����|4�[�����:�e�n�u�w�-�@�������WF��~ ��!�����n�u�w�-�@��Cӯ��`2��{!��6�����u�d�w�2����I��ƹF��hY��*���#�1�o��w�	�(���0��ƹF��hY��U���������!���6���F��@ ��U���_�u�u�
����������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��V�����u������4�ԜY�Ƽ�9��T��;ʆ�������8���H�ƨ�D��^����u�
�
�e�6�����Y����g"��x)��N���u�%�b�d�w�}�9ύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����W��G1�����u��
���L���YӖ��lW��N��U���
���
��	�%���Lӂ��]��G�U���%�b�d�
�'�+���0�Ɵ�w9��p'�����u�
�
�f�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ѓ� 9��h��U���������}���Y����R�'��&���������W��Y����G	�UךU���
�
�a�4��1�W���7ӵ��l*��~-�U���%�b�d�u�w��$���5����l0��c!��]���1�"�!�u�~�W�W���&Ĺ��l��A��Oʜ�u��
���f�W���	���)��=��*����n�u�u�'�e��������|3��d:��9����_�u�u��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�
9��h��U���������}���Y����\��b:��!�����
����_������\F��d��Uʥ�d�
�%�#�3�g�8���*����|!��d��Uʥ�d�u�u����;���:����g)��_����!�u�|�_�w�}�(�������WF��~ ��!�����n�u�w�-�F���Y����g"��x)��N���u�%�d�
�'�+���0�Ɵ�w9��p'�����u�
�`�o��	�$���5����l0��c!��]���1�"�!�u�~�W�W���&�ӓ�C9��SN�:��������t�}���B����A��C�� ���7�=�#�:�w�h�6���@������=N��U���'�7�!�u���0���+����}9��q!��U�����_�u�w�)�����Ə�a#��r ��4������u�1�?����CӇ��[��T��ʼ�_�u�u�8��d�6֝�&�ʤ�@9��h\�@��.��
����.�������5��y>��*����h�y����"���0����J��d1��%�����h�6�-�o����A����{*��~ ��!�����g�{�g�m�GÖ�*����f2��e-�����'�y��
���;���D����
V��&��*���
��h�b���$���-����\��"��&�����e����9���)����5��n ��3��b������#��@���9F������!�4�
�:�$�����&����`2��{!��6��u�d�n�u�w�>�����ƭ�l��D�����
�u�u����>���D����l�N�����;�u�%���)�(���&����`2��{!��6�����u�d�3�*����P���V��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�l��������\�_�N���u�6�;�!�9�}��������EU��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��h_��U���
���
��	�%���Y����G	�N�U��n�u�u�6�9�)����	����@��A_��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�F��Cӵ��l*��~-��0����}�u�:�9�2�G���D����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����L���5��h"��<������}�w�2����I����D��^�N���u�6�;�!�9�}��������ER��T��!�����
����_�������V�S��E��w�_�u�u�8�.��������]��[��D��������4���Y����\��XN�U��w�e�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�f��}���Y����G�������!�9�a�f�m��3���>����v%��eN��U���;�:�e�u�j��G��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���f�1�"�!�w�t�M���I����l�N�����;�u�%�6�9�)����L����g"��x)��*�����}�u�8�3���Y���W��UךU���:�&�4�!�6�����&����F��d:��9�������w�n��������\�^�E��u�u�6�;�#�3�W�������l
��hY��U���
���
��	�%���Y����G	�N�U��d�w�_�u�w�2����Ӈ��P	��C1��A��o������!���6�����Y��E���h�w�e�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�f�m�U�ԜY�Ư�]��Y�����;�!�9�a��g�$���5����l0��c!��]���:�;�:�e�w�`�U��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�f�1�"�#�}�^��Y����D��N�����!�;�u�%�4�3����M���5��h"��<������}�w�2����I����D��^�����u�:�&�4�#�<�(���
����9��N��1��������}�DϺ�����O�
N��D��n�u�u�6�9�)����	����@��AZ��U����
�����#���Q�ƨ�D��^��O���d�d�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������pF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��rN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��_�E��u�u�6�;�#�3�W�������l
��1��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�D��n�u�u�6�9�)����	����@��A[��E��������4���Y����\��XN�U��w�e�e�w�]�}�W���
������T�����`�d�o����0���/����aF�
�����e�u�h�w�g�m�U�ԶY����Z��[N��*���3�8�o����0���/����aF�
�����e�u�h�w�f�f�W�������Q����*���:�<�2�o�$�/���Y����G��U��U���
�;�:�<�0�2�W���:����^F��D�����&�w�:�0�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����A����|)��v �U���&�2�4�u���(���
���5��h"��<������}�b�9� ���Y����F�D�����
�
�
�'�0�g�$���5����l0��c!��]���1�"�!�u�~�g�W��I����V��^�E��u�u�&�2�6�}�(߁�&����_��Y1���������W�W���������h^�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
����������g"��x)��*�����}�`�3�*����P���F��P ��U���
�
�'�2�m��3���>����v%��eN��@ʱ�"�!�u�|�m�}�G��I����V��^�N���u�&�2�4�w��(ށ�	����l��D��Oʆ�����]�}�W�������lV��h�����%�0�u�u���8���Y���A��N�����4�u�
�
��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*ڊ�
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u���(�������]9��PN�&������_�w�}����Ӗ��lT��G1�����0�u�u����>���D����l�N�����u�
�
�
�9�.���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T����*ي�'�2�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��d��Uʦ�2�4�u�
����������@��N��1�����_�u�w�4����	�֓�l��A�����u�u��
���W��^����F�D�����
�
�
�;�$�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��h^��*���2�o�����4���:����W��S�����|�o�u�e�g�m�G��I����D��N�����4�u�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�I�ғ�C9��S1�����u��
���}�J���^���F��P ��U���
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h[�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1����L����E
��G��U����
���w�`�P���s���@��V��*ڊ�
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lV��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*݊�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��lQ��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�m�@���&����C��T��!�����u�h�p�z�}���Y����R
��h^��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�֓�l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G���s���@��V��*ڊ�
�%�#�1�>�����Y����)��tUךU���<�;�9�%�g�e��������V�=��*����u�h�r�p�W�W���������hW�����2�o�����4���:����W��S�����|�_�u�u�>�3�Ϯ�I�ߓ�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*ӊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�e�n�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lV��1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&�֓�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*���4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
��m��������V�=��*����u�h�r�p�W�W���������h_�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ù��l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G���s���@��V��*ڊ�d�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���F���&����C��T��!�����u�h�p�z�}���Y����R
��h^��G���
�<�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����T��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�g�4�
�;���������g"��x)��N���u�&�2�4�w��(�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�f�4��1�(���
���5��h"��<��u�u�&�2�6�}�(߁�J����E
��G��U����
���w�`�P���s���@��V��*ڊ�a�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��Z�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�a�6���������\��c*��:���n�u�u�&�0�<�W���&�ғ�C9��S1�����u��
���}�J���^���F��P ��U���
�`�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�*���2�o�����4���:����W��S�����|�o�u�e�g�m�G��I����D��N�����4�u�
�
�b�<�(���&����Z�=��*����n�u�u�$�:����&ù��l��A�����u�u��
���W��^����F�D�����
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�l��������V�=��*����u�h�r�p�W�W���������h^�����2�o�����4���:����W��S�����|�_�u�u�>�3�Ϯ�L�֓�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*ڊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�`�g�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lS��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����H����TF��d:��9�������w�l�W������F��L�E��e�e�e�e�g��}���Y����R
��h[��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�`�d�6��������5��h"��<���h�r�r�_�w�}����Ӗ��lT��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�B���	����	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�u�W�W���������h\�����1�<�
�<�w�}�#���6����9F������%�`�g�4��1�(�������g"��x)��U��r�r�_�u�w�4����	�ӓ�l��D��Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�h�D�������`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�w�]�}�W�������lS��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�`�f�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L�ғ�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�b�i����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��lR��G1�����
�<�u�u���8���B�����Y�����a�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����L����@��N��1��������}�F�������V�=N��U���;�9�%�`�b�-����Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�w�_�u�w�4����	�ӓ�l��A�����<�u�u����>��Y����Z��[N��@���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�B�������TF��d:��9�������w�l�W������]ǻN�����9�%�`�c�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�L�Г�C9��S1��*���u�u��
���L���Yӕ��]��G1��C���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�h�@���&����	F��s1��2������u�f�}�������9F������%�`�b�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����N����E
��^ �����u��
���f�W���
����_F��1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�b�e��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�`�m�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�B�������W9��h��U����
���l�}�Wϭ�����C9��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�`�n�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����l�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�h�N���&����Z��^	��U���
���n�w�}�����Ƽ�9��V�����'�2�o����0���C���]ǻN�����9�%�`�d��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*ߊ�e�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�h�F߁�	����l��D��Oʆ�����]�}�W�������lS��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�`�f���������g"��x)��*�����}�`�3�*����P���F��P ��U���
�d�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�B��&����_��Y1���������W�W���������h_�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�b�l�(���
���5��h"��<������}�b�9� ���Y����F�D�����
�
�g�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����H����l��h�����o������}���Y����R
��h[��G���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�h�F܁�����\��c*��:���
�����h��������l�N�����u�
�
�f�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�L����R��[
�����2�o�����4�ԜY�ƿ�T����*���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�B��&����Z�=��*����
����u�BϺ�����O��N�����4�u�
�
�c�-����Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�w�_�u�w�4����	�ӓ�9��h��*���&�2�o����0���s���@��V��*ߊ�a�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����Hƹ��l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��h����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��lW��V�����;�&�2�o���;���:���F��P ��U���
�`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N�֓�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�`�m����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��lV��G1�����
�<�u�u���8���B�����Y�����e�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����H����@��N��1��������}�F�������V�=N��U���;�9�%�b�f�-����Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�w�_�u�w�4����	�ѓ�l��A�����<�u�u����>��Y����Z��[N��B���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�@�������TF��d:��9�������w�l�W������]ǻN�����9�%�b�g�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�N�ԓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��G���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�j�D���&����	F��s1��2������u�f�}�������9F������%�b�f�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����J����E
��^ �����u��
���f�W���
����_F�� 1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�`�i��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�b�a�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�@�������W9��h��U����
���l�}�Wϭ�����C9��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�b�b�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����`�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�j�B���&����Z��^	��U���
���n�w�}�����Ƽ�9��V�����'�2�o����0���C���]ǻN�����9�%�b�c�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��B���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�`�k��������l��T��!�����n�u�w�.����Y����9��h��*���2�o�����4��Y���9F������%�b�b�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��B���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b�`�<�(���&����Z�=��*����n�u�u�$�:����&Ĺ��R��[
�����o������M���I��ƹF��^	��ʥ�b�m�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F�� 1�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�b�m�6���������\��c*��:���n�u�u�&�0�<�W���&˹��l��h���������g�W��B�����Y�����l�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b�l�4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�&����_��E��Oʆ�����m�}�G��Y����Z��[N��B��
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lQ��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b�d�
�'�+����&����	F��s1��2���_�u�u�<�9�1����Hù��l��h���������g�W��B�����Y�����d�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h_�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�b�d��-��������TF��d:��9����_�u�u�>�3�Ϯ�N����R��[
�����o������M���I��ƹF��^	��ʥ�b�d�
�;�$�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��hY��G���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b�f���������@��N��1�����_�u�w�4����	�ѓ�9��h��*���2�o�����4��Y���9F������%�b�d�
�9�.���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T����*���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�`�l�(�������]9��PN�&������_�w�}����Ӗ��lW��V�����'�2�o����0���C���]ǻN�����9�%�b�d��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*݊�a�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�j�Fہ�	����l��D��Oʆ�����]�}�W�������lQ��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�b�f���������g"��x)��*�����}�`�3�*����P���F��P ��U���
�`�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�@��&����_��Y1���������W�W���������h_�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�n�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�n�<�(���&����Z�=��*����n�u�u�$�:����&ʹ��l��h���������g�W��B�����Y����
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lW��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�l�(�������A��N��1�����o�u�g�f�W���
����_F��\�����2�o�����4�ԜY�ƿ�T����G���0�u�u����>���D����l�N�����u�
�g�4��1�(���
���5��h"��<��u�u�&�2�6�}�(�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����������:�#�(�(���I����g"��x)��*�����}�u�8�3���Y���D��N�����4�u�%�&�0�?���M����|)��v �U���&�2�4�u�%���������lS��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:��������\
��E!��*���e�'�2�g�`�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h������!�`�
��8�(��A����g"��x)��*�����}�u�8�3���B�����Y�����7�:��'�"��D�������^��N��1��������}�GϺ�����O��N�����4�u�'�
�8�1�������� 9��P1�M���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<��������|��]��*���
�e�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����Q	��v�� ���f�`�'�2�e�d�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����'��!�`������H���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�7�:��%�(�(���N����lT��N�&���������W������\F��d��Uʦ�2�4�u�'��2����6���� 9��E��G��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������A��C1�*ӊ�0�
�d�m�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��X�����
�f�d�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����:��'� ��n�Fށ�����^�=��*����
����u�W������]ǻN�����9�4�'�7�8�����&�Փ�9��P1�F���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<��������|��]��F���2�g�f�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��[/��:���`�
�a�'�0�o�C���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���9�'��!�b��B�������F��d:��9�������w�m��������l�N�����u�'�
�:�;�/�8���L¹��U��X��D��������4���Y����\��XN�N���u�&�2�4�w�/�(�������F��1�����g�`�u�u���8���&����|4�N�����u�|�_�u�w�4��������\	��E�����
�
�0�
�f�e�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1�����'� �
�d�e�/���O����`2��{!��6�����u�e�3�*����P���F��P ��U���
�:�9�'��)�Bށ�&����W��T��!�����
����_�������V�=N��U���;�9�4�'�5�2�6�������lR��R	��D��o������!���6�����Y��E��u�u�&�2�6�}��������A)��h[��@���2�g�b�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��[/��:���`�
�
�0��l�D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V������'� �
�f�j����K����	F��s1��2������u�g�9� ���Y����F�D�����'�
�:�9�%����&˹��T9��]��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�?��������W��h��*��m�o�����4���:����V��X����n�u�u�&�0�<�W���&����r��B��D��
�0�
�g�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��U��4��� �
�d�d��8�(��A����g"��x)��*�����}�u�8�3���B�����Y�����7�:��'�"��F��&����T��T��!�����
����_�������V�=N��U���;�9�4�'�5�2�6�������lW��E��G��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������A��C1�*���'�2�g�g�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��X�����!�`�
�`�%�:�E��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����:�9�'��#�i�(߁�����l��N��1��������}�GϺ�����O��N�����4�u�'�
�8�1��������9��P1�F���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<��������|��W��*���
�g�m�o���;���:����g)��^�����:�e�n�u�w�.����Y����Q	��v�� ���l�g�'�2�e�i�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����'��!�a������K���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�7�:��%�(�(���M����lT��N�&���������W������\F��d��Uʦ�2�4�u�'��2����6����
9��E��G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������A��C1�*܊�0�
�g�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��X�����
�l�b�'�0�o�A���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���9�'��!�c��(���&����\��c*��:���
�����}�������9F������4�'�7�:��/����@�ߓ�V��Y�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%���������lR��^�����g�f�o����0���/����aF�
�����e�n�u�u�$�:��������\
��E!��*���d�
�0�
�e�e�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1�����'� �
�l�f�����K���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�7�:��%�(�(���H����T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�?��������_��1����e�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����_'��x��Aӊ�`�'�2�g�g�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������[�����:�%�d�
�"�l�E߁�K����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���݁�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������l ��h"�����'�2�c�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʃ�Z��Y
�����d�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��9��V
�����3�
�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��[�����:�%�g�
�b�;�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����!��'��8��@�������P��N�&���������W������\F��d��Uʦ�2�4�u�8��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�9�
�:��2���&�ӓ�l ��]�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%���������C9��h_��G���
�a�u�u���8���&����|4�N�����u�|�_�u�w�4��������G9��E1�����b�d�
�
�"�o�C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��B�������F��d:��9�������w�m��������l�N�����u�'�
�!��/�;���&�ѓ�9��Q��@���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��Dߊ�
� �g�c�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�g�
�`�`�;�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����!��'��8��@��&˹��lT��T��!�����
����_�������V�=N��U���;�9�4�'�;���������9��hW�� ��m�o�����4���:����V��X����n�u�u�&�0�<�W���&����\��X��G݊�`�d�
� �e�o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g��h�Fށ�����\��c*��:���
�����}�������9F������4�'�9�
�8�����KĹ��lW��Q��M���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<����&����	��h\��Dߊ�f�3�
�m�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��C1�����:�
�b�d��i����A����`2��{!��6�����u�e�3�*����P���F��P ��U���
�!��'��2�(���Hƹ��l ��W�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%���������C9��h_�����l�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����u	��{��*���e�3�
�g�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�l�(ށ�����\��c*��:���
�����}�������9F������4�'�9�
�8�����Kʹ��lT��B1�A��������4���Y����\��XN�N���u�&�2�4�w�/�(���?����\	��W��@���3�
�e�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l
��q��9���
�l�d�
��(�D��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�:�
�:�'�o�(���L���� W��N��1��������}�GϺ�����O��N�����4�u�'�
�#���������lW��1��*��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������A9��X��L��
�
� �f�c�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��[�����:�%�g�
�b�e����K����`2��{!��6�����u�e�3�*����P���F��P ��U���
�!��'��2�(���Hƹ��U��\��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�1�(���&����lT��[��E���
�f�u�u���8���&����|4�N�����u�|�_�u�w�4��������G9��E1�����l�d�
�d�1��C���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*����'��:��d�Fځ�K���� R��N��1��������}�GϺ�����O��N�����4�u�'�
�#���������lW��]�� ��m�o�����4���:����V��X����n�u�u�&�0�<�W���&����\��X��Gӊ�`�d�
� �d�o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g��h�Fځ�����\��c*��:���
�����}�������9F������%��&�9���(���H����CW��N��1��������}�F�������V�=N��U���;�9�%��$�1�(ف�&����_��G_�Oʆ�������8���H�ƨ�D��^����u�<�;�9�5�2�(��� ����Q��B1�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����|��Y�����3�
�f�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q	��h�����
�b�3�
�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��B9��0���� �
�l�1��B߁�J����g"��x)��*�����}�`�3�*����P���F��P ��U���
�:�9�'��)�Cց�����l ��[�����u��
����2���+������Y��E��u�u�&�2�6�}� ���&����	��h_�����d�e�%�m�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������d9��h(��*���%�d�
� �f�h�(��Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����!��'��8��G���&����l��T��!�����
����_������\F��d��Uʦ�2�4�u�:�;�%�#�������U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?��������l*��G1�*���d�l�
�d�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������\	��O"��:���a�
� �d�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��*����'��:��i����K�ޓ�^�=��*����
����u�W������]ǻN�����9�7�:�
�8�8����&�ғ�F9�� Z��G��������4���Y����\��XN�N���u�&�2�4�w�2����&����	��h\�����g�e�%�m�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�\
��X
�����
�b�3�
�e�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*��� �d�g�
�e�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������y=�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�<�(���&����W��N��:����_�u�u�>�3�Ͽ�&����Q��Z�U������n�w�}�����ƭ�l��h��*��o�����W�W���������D�����m�l�o����9�ԜY�ƿ�T�������7�1�d�b�m��8���7���F��P ��U���&�2�7�1�f�k�MϜ�6����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w�-��������U�,��9���n�u�u�&�0�<�W���
����W�� \��U�����n�u�w�.����Y����Z��S
��C������]�}�W�������C9��P1�����u�u����f�W���
����_F��h��*���
�a�o����9�ԜY�ƿ�T�������7�1�b�u�w��;���B�����Y�����<�
�1�
�e�g�5���<����F�D�����%�&�2�7�3�d�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����W��N��:����_�u�u�>�3�Ͽ�&����Q��W�Oʗ����_�w�}����Ӈ��@��U
��@��o�����W�W���������D�����d�d�o����9�ԜY�ƿ�T�������7�1�d�e�m��8���7���F��P ��U���&�2�7�1�e�m�MϜ�6����l�N�����u�%�&�2�5�9�E��CӤ��#��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-��������Q�,��9���n�u�u�&�0�<�W���
����W��X��U�����n�u�w�.����Y����Z��S
��G���u����l�}�Wϭ�����R��^	�����l�u�u����L���Yӕ��]��V�����1�
�e�u�w��;���B�����Y�����<�
�1�
�f�}�W���5����9F������4�
�<�
�3��E���Y����v'��=N��U���;�9�4�
�>�����J����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�G������]�}�W�������C9��P1����d�o�����}���Y����R
��G1�����1�f�a�o���2���s���@��V�����2�7�1�a�c�g�5���<����F�D�����%�&�2�7�3�i�D��;����r(��N�����4�u�%�&�0�?���K����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lR��T��:����n�u�u�$�:����	����l��hZ�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�`�u�u���6��Y����Z��[N��*���
�1�
�c�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��j�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&���� _��N��:����_�u�u�>�3�Ͽ�&����Q��^�Oʗ����_�w�}����Ӈ��@��U
��A���o�����W�W���������D�����a�e�o����9�ԶY����\��Y��U����l�l�3�g�0����ד�V
��X��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�l� ���1����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�<�f����Mϗ�-����l�N��Uʱ�;�
���w�}�9���<��ƹF�N��������o��	�0���s���F�S��*����u�u����L���Y����� 1��1���o�����W�W���Y�ƨ�]^��~*��U������n�w�}�W�������d/��N�<�����_�u�w�}�W���Hù��w2��N��!����_�u�u�w�}���&����{F��~ ��2���_�u�u�u�w�4�F݁�0����	F��c+��'�ߊu�u�u�u�>�l�(���-����z(��p+�����u�u�u�<�f��>���Y�ƅ�g#��eUךU���u�u�<�d���#���Y����t#��=N��U���u�<�d�
��	�W���7����a]ǻN��U���<�d�
���}�W���<����9F�N��U���!����m��#���+����F�G��U�ߊu�u�u�u�>�l�Mϗ�Y����)��t1��6���u�d�u�:�9�2�G��Y���F��^ �Oʜ�u��
����2���+������Y��E��u�u�u�u�3�3�W���7ӵ��l*��~-��0����}�`�1� �)�W���s���F�S��U���������!���6���F��@ ��U���_�u�u�u�w�4�B��0�Ɵ�w9��p'��#����u�d�u�8�3���B���F�
��C���u��
���(���-���S��X����n�u�u�u�w�9����Y����g"��x)��*�����}�`�3�*����P���F�N�����u������4���:����W��S�����|�_�u�u�w�}���Cӯ��`2��{!��6�����u�d�w�2����I��ƹF�N����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���H����z(��c*��:���
�����h��������l�N��Uʱ�;�g�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������\��yN��1��������}�F�������V�=N��U���u�<�d�u�w��$���5����l0��c!��]���1�"�!�u�~�W�W���Y�ƨ�]W��N��U���
���
��	�%���Lӂ��]��G�U���u�u�1�;�a�g�>���-����t/��a+��:���d�u�:�;�8�m�L���Y�����Y��U���������4���Y����\��XN�N���u�u�u�1�"�}�W���Y����)��t1��6���u�d�u�:�9�2�G���B����������;�n�_�u�w�>��������'��/�����8�-�d�!�f�.�ہ�&�ƅ�9F�	�����u�_�u�u�w�}�3��0����v4��N��U��������g�>���>����F�N�����
���u�w��2���B���F�
��G�����o����%�ԜY���F��Y]��<���u�u����f�W���Y����Z��`'��=������]�}�W���Y����l1��c&��U�����n�u�w�}�WϺ�Ź��w2��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�n�
�3���Cӯ��v!��d��U���u�1�;�e� ��?��0����v4��N��U���1�;�d����Mϗ�-����l�N��Uʱ�;�g����g�>���>����F�N�����f����m��#���+���F�N��������o��	�0���s���F�S��@�����o����%�ԜY���F��Y_��"����o�����}���Y���W�� 1��1���o�����W�W���Y�ƨ�F��~*��U������u�l�}�WϮ����F�N�����u�u�����0���/����aF�
�����e�n�u�u�w�}����Y�ƅ�5��h"��<������}�w�2����I��ƹF�N����o��u����>���<����N��S�����|�_�u�u�w�}���Cӯ��`2��{!��6�����u�e�3�*����P���F�N�����u������4���:����V��X����n�u�u�u�w�9����Y����g"��x)��*�����}�u�8�3���B���F�
��B���u��
���(���-���F��@ ��U���_�u�u�u�w�4�O��0�Ɵ�w9��p'��#����u�e�1� �)�W���s���F�S��U���������!���6�����Y��E��u�u�u�u�3�3�G��0�Ɵ�w9��p'��#����u�e�1� �)�W���s���F�S��D���u��
���(���-���F��@ ��U���_�u�u�u�w�4�F���Y����g"��x)��*�����}�u�8�3���B���F�
��D���u������4���:����V��X����n�u�u�u�w�9���Cӯ��`2��{!��6�����u�e�3�*����P���F�N�����o��u����>���<����N��S�����|�_�u�u�w�}���Y�ƅ�5��h"��<������}�w�2����I��ƹF�N����u�u�����0���/����aF�
�����e�n�u�u�w�}����Y�ƃ�gF��s1��2������u�g�9� ���Y���l�N��ʶ�8�:�0�!�]�W������� ��h��*���:�
�0�a�f��(��CӅ��C	��Y��@���l�l�3�e�:�%�F٪�H����9��h_ךU���0�0�<�u�6�}�}���Y���z"�	N����u�u�u� ��	�0���G����F�N�����
���u�i�l�[���Y�����1��1���h�u�c�_�w�}�W����Փ�z"��S�D���u�u�u�u�3�3�(���-���W��=N��U���u�<�`����J���O���F�N��܊���u�k�f�q�W���Y����Z��`'��=��u�c�_�u�w�}�W���A����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���<�d�
���}�I��U���F�
��Dۊ���u�k�f�q�W���Y����Z��h9��!���k�d�y�u�w�}�WϺ��Փ�z"��S�D���u�u�u�u�3�3�C���=���F��d��U���u�1�;�`� ��?��Y����F�N�����c����j�}�A�ԜY���F��Y_��"����h�u�y�w�}�W�������d/��N��U��_�u�u�:�#�0����Y���F��^ �H���
�
�
�;�$�:�}���Y���W��S����d�<�
�<�{�}�W���Yӂ�� F���*؊�;�&�2�_�w�}�W������F��1�����<�y�u�u�w�}����Y����lV��h�����_�u�u�u�w�4�A��Y����9��h��Y���u�u�u�1�9�}�IϮ�I�Г�]9��PBךU���u�u�<�m�j�}�(߁�&����Z�N��U���1�;�u�k�'�m�O���&����9F�N��U���d�u�k�%�g�d������ƹF�N����u�k�%�e�f��������F�N����h�u�
�
�f�4�(���U���F�
��D���k�%�e�d��3����s���F�S��A��u�
�
�f�>����Y���F��^ �U��%�e�d�
�9�.��ԜY���F��Y_�H���
�
�`�<��4�[���Y�����Y��Kʡ�%�3�
�d�a�-�[���Y�����CN��U���9�
�:�
�8�-�Fف�����9��G����u�
�
� ��k�ށ��ғ�9��b_��U���%�;�;�u�b��N����֓�F����*���a�d�
�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���W��=N��U���u�<�g����J���O���F�N��ي���u�k�f�q�W���Y����Z��`'��=��u�c�_�u�w�}�W���L����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���<�b����`�W��s���F�S��*����u�k�d�{�}�W���Yӂ��
9��s:��H���c�_�u�u�w�}���&����{F�_����u�u�u�<�f��>���Y���JǻN��U���<�d�
���}�I��U���F�
��Dي���u�k�f�q�W���Y����Z��h9��!���k�d�y�u�w�}�WϺ��ӓ�z"��S�D���u�u�u�u�3�3�A���=���F��d��U���u�1�;�b� ��?��Y��ƹF�N��������h�w�k�}���Y������FךU���u�u�<�d�j�}�(ځ�&����Z�N��U���1�;�u�k�'�h�F���&����9F�N��U���f�h�u�
���������F�N�����k�%�`�f�>����Y���F��^ �H���
�
�
�;�$�:�}���Y���W��S����`�<�
�<�{�}�W���Yӂ��F���*܊�;�&�2�_�w�}�W������F��1�����<�y�u�u�w�}����Y����lS��h�����_�u�u�u�w�4�F���GӖ��l_��Y1���ߊu�u�u�u�>�l�W���	�ӓ�9��h��Y���u�u�u�1�9�o�J���&ƹ��l��D�����u�u�u�<�f�}�IϮ�L����Z��^	�U���u�u�1�;�c�`�W���&�Փ�]9��PBךU���u�u�<�d�w�c����Hǹ��l��d��U���u�1�;�c�j�}�(ځ�L����@��=N��U���u�<�d�u�i�)����&����l��=N��U���u�:�!�h�w�
��������\��1��*��g�%�m�n�]�}�W���&����P��1��ފ�c�d� �u�w�2�����ơ�r'��vW��*ڊ� �
�c�:��8�C��&���F��Y��ʸ�%�}�u�u�w�}�>���G����F�N��;������h�w�q�W���Y����Z��`'��=��u�c�_�u�w�}�W���K����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���<�a����`�W��s���F�S��*����u�k�d�{�}�W���Yӂ��9��s:��H���c�_�u�u�w�}����.����[�X�U���u�u�1�;���#���G����9F�N��U���l����j�}�A�ԜY���F��Y_��"����h�u�c�]�}�W���Y����9��s:��H���c�_�u�u�w�}���&����{F�_����u�u�u�<�f��>���Y���JǻN��U���<�d�
���}�I��U���F�
��Dߊ���u�k�f�q�W���Y����Z��h9��!���k�d�y�u�w�}�WϺ��ѓ�z"��S�A�ߊu�u�u�u�8�)� ���1���P�N�����u�4�u�_�w�}�W������F�� 1�����<�y�u�u�w�}����Y����lQ��h�����_�u�u�u�w�4�D��Y����9��h��Y���u�u�u�1�9�}�IϮ�N�Փ�]9��PBךU���u�u�<�`�j�}�(؁�&����Z�N��U���1�;�u�k�'�j�B���&����9F�N��U���b�h�u�
���������F�N�����k�%�b�b�>����Y���F��^ �H���
�
�
�;�$�:�}���Y���W��N��U���
�
�;�&�0�W�W���Y�ƨ�]W��
P��*݊�e�<�
�<�{�}�W���Yӂ��T�	N��B��
�;�&�2�]�}�W���Y���� F���*���<�
�<�y�w�}�W�������[�G1��Dي�;�&�2�_�w�}�W�������X��hY��A���
�<�y�u�w�}�WϺ����F�� 1�*���&�2�_�u�w�}�W���H�����h��D��
�d�_�u�w�}�W������Z1��C1�����:�
�e�3��l�C���A��ƓF�Q1�����d�!�d�&�;��(ށ�J����\��Y��U����l�l�3�g�0����ד�V
��1�U���2�;�'�6�:�-�_���Y���/��
P��Y���u�u�u����6���D����9F�N��U���d����j�}�[���Y�����1��1���h�u�y�u�w�}�WϺ�����w2��
P��Y���u�u�u�1�9��>���Y���l�N��Uʱ�;�
���w�c�F�ԜY���F��YX��<���u�k�d�_�w�}�W����ѓ�z"��S�D�ߊu�u�u�u�>�e� ���1���JǻN��U���<�l����`�W��Y���F��^ �*����u�k�d�]�}�W���Y����9��s:��H���y�u�u�u�w�9����.����[�BךU���u�u�<�d���#���G����F�N�����a����j�}�[���Y�����[��<���u�k�d�_�w�}�W�������d/��N��U���u�u�u�u�3�3�@���=���F��=N��U���u�:�!����J���P�����CN�����u�u�u�u�3�3�W�������\	��E����
�
�0�
�e�n�}���Y���W��S����7�:��'�"��N�������U��=N��U���u�<�f�h�w�/�(�������F��1�����g�a�y�u�w�}�WϺ������h������!�a�
��8�(��A���F�N�����k�4�'�7�8�����&�ߓ�l��h\�F�ߊu�u�u�u�>�k�J�������\
��E!��*���`�'�2�g�b�q�W���Y����Z��
P�����:�9�'��#�i�(ف�����U�N��U���1�;�u�k�6�/����8����G9��hY�����g�m�_�u�w�}�W���@���R��U��4��� �
�l�m�%�:�E��U���F�
��D���k�4�'�7�8�����&�ߓ�l��h\�M�ߊu�u�u�u�>�l�W�������\	��E����
�e�'�2�e�e�[���Y�����\��Kʴ�'�7�:��%�(�(���H¹��T9��V�U���u�u�1�;�d�`�W���&����r��B��L��
�0�
�g�d�W�W���Y�ƨ�]W��
P�����:�9�'��#�i�(�������_��=N��U���u�<�d�u�i�<��������|��W��A���2�g�e�y�w�}�W�������[�V������'� �
�n�l�(���&����l�N��Uʱ�;�b�h�u�:����KŹ��l�N��Uʱ� �u�k�7�8���������C9��h��D��
�d�|�_�w�}����������h��A���d� �u�u�8�-����Y�Ӎ�
_��t��*���
�c�:�
�2�i�F��Y����V��^�����_�u�u�u�w��J���U���F� ��*����u�k�d�]�}�W���Y����l1��c&��K��_�u�u�u�w�4�E���=���F��=N��U���u�<�f����J���U���F�
��A�����h�u�{�}�W���Yӂ��9��s:��H���y�u�u�u�w�9�ف�0����X�d��U���u�1�;�
��	�W���H���F�N��Ҋ���u�k�f�W�W���Y�ƨ�]_��~*��U��d�_�u�u�w�}���&����{F�_�U���u�u�1�;�f�
�3���D����9F�N��U���d�
���w�c�F�ԜY���F��Y_��"����h�u�y�w�}�W�������l1��c&��K��_�u�u�u�w�4�Fځ�0����X�d��U���u�1�;�c� ��?��Y��ƹF�N����
���u�i�i�}���Y���W	��h9��!���k�d�_�u�w�2�ϳ�	��ƹF�N����h�u�'�
�8�1��������9��P1�@���u�u�u�u�3�3�W�������\	��E�����
�
�0�
�f�e�}���Y���W��S����7�:��'�"��F�������P��=N��U���u�<�a�h�w�/�(�������F��1�����g�c�y�u�w�}�WϺ������h������!�`�
��8�(��J���F�N�����k�4�'�7�8�����&�ד�l��h\�M�ߊu�u�u�u�>�j�J�������\
��E!��*���c�'�2�g�o�q�W���Y����Z��
P�����:�9�'��#�h�(؁�����^�N��U���1�;�u�k�6�/����8����G9��hV�����d�f�_�u�w�}�W���H�����h������!�`�
��8�(��A���F�N����h�u�'�
�8�1��������V��R	��G��_�u�u�u�w�4�F���GӇ��l��[/��:���`�
�d�'�0�o�G��Y���F��^ �U��4�'�7�:��/����H����A��\�Y���u�u�u�1�9�i�J�������\
��E!��*���d�
�0�
�e�e�}���Y���W��N��U���
�:�9�'��)�Bށ�M����lT��BךU���u�u�<�d�w�c��������A��C1�*���'�2�g�g�{�}�W���Yӂ��Q�	N�����
�d�c�%�{�}�W���Yӂ��GF������
�:�
�:�'�o�(���H����CW��dךU���
�
� �
�a�2�(���M�ד�l3��N�����0�!�8��n��4���&����P��1��ފ�
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�_�U���u�u�1�;���#���G����F�N�����
���u�i�l�}���Y���W��h9��!���k�d�_�u�w�}�W���M����g.�	N����u�u�u�<�b�
�3���D����9F�N��U���c����j�}�[���Y����� 1��1���h�u�y�u�w�}�WϺ�˹��w2��
P��Y���u�u�u�1�9��>���Y���l�N��Uʱ�;�e����`�W��Y���F��^ �*����u�k�d�]�}�W���Y����9��s:��H���y�u�u�u�w�9����.����[�BךU���u�u�<�d���#���G����F�N�����`����j�}�[���Y�����X��<���u�k�d�_�w�}�W�������d/��N��U���u�u�u�u�3�(�(���-���W�N�����u�4�u�_�w�}�W������F��E1�����'� �
�f�g�/���N��ƹF�N����h�u�'�
�8�1��������9��P1�B���u�u�u�u�3�3�W�������\	��E�����
�
�0�
�g�n�}���Y���W��S����7�:��'�"��D�������^��=N��U���u�<�`�h�w�/�(�������F��1�����g�l�y�u�w�}�WϺ������h������!�`�
��8�(��A���F�N�����k�4�'�7�8�����&�Փ�l��h\�F�ߊu�u�u�u�>�e�J�������\
��E!��*���b�'�2�g�g�q�W���Y����Z��
P�����:�9�'��#�h�(ׁ�����U�N��U���1�;�e�h�w�/�(�������F��1�����g�d�y�u�w�}�WϺ����F��E1�����'� �
�f�f�����H����F�N�����g�h�u�'��2����6���� 9��h��*��m�_�u�u�w�}���Y����A��X�����!�`�
�g�%�:�E��U���F�
��D���k�4�'�7�8�����&�Փ� 9��P1�F���u�u�u�u�3�3�B��Y����Q	��v�� ���f�d�
�0��l�D�ԜY���F��Y_�H���'�
�:�9�%����&�ӓ�V��Z����u�u�u�<�f�}�IϪ�	����W��h����u�u�u�:�#�`�W�������u	��{��*���3�
�g�e�'�e�L�Զs���F���U���'�;�u�!�#�}����*����F����U���!�u�4�=�9�s�Z�ԜY�ƭ�l%��Q�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�u�u�w�}�W���Y���F���6���&�u�h�4������s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������TF��D��U���6�&�{�x�]�}�W���&ù��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g�m��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lV��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����lV��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����9��R	�����;�%�:�0�$�}�Z���YӖ��lV��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�e�g�-����DӇ��P	��C1��D܊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�G1��E���
�9�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\���!�0�u�u�w�}�W���Y���F���*ڊ�'�2�i�u���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�d��-����	����R��P �����&�{�x�_�w�}�(߁�I����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��m��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lV��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����g�|�!�0�w�}�W���Y���F�N��U���u�
�
�e�6��������F��1�*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��^�����4�&�2�u�%�>���T���F��1�*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G��&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h^��E���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�e�'�8�W��	�֓�]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����H¹��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��_�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Q����Z��S
��F���!�0�u�u�w�}�W���Y���F�N��U���
�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�H����E
��G��U��%�e�d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e�d�
�'�0�<����Y����V��C�U���%�e�d�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�d�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(߁�H����TF���*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h_�����9�
�'�2�6�.��������@H�d��Uʥ�e�d�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��D؊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F��*���
�1�
�f�~�)����Y���F�N��U���u�u�u�u���E���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9��\�����1�%�0�u�j�-�G��&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�F݁�����@��YN�����&�u�x�u�w�-�G��&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�g�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(߁�K����E
��G�����_�u�u�u�w�}�W���Y���C9��\�����i�u�
�
�e�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�f�4��1�(���Ӈ��Z��G�����u�x�u�u�'�m�F܁�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�e�d��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����J����[��=N��U���u�u�u�u�w�}�W���Y����U��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��Uʥ�e�d�
�%�!�9����Y����lV��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lW��G��U���<�;�%�:�2�.�W��Y����lV��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���D��������T�����d�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��]�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e�d�
�'�0�a�W���&����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������W9��R	�����;�%�:�0�$�}�Z���YӖ��lW��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����Hǹ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�Wǿ�&����Q��]�U���;�_�u�u�w�}�W���Y���F�N��E��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�d�d�}����s���F�N��U���u�u�u�u�'�m�Fہ�	����l��PN�U���
�a�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ڊ�a�%�0�u�$�4�Ϯ�����F�=N��U���
�a�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����R��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�e�d�
�%�!�9�^������F�N��U���u�u�u�u�'�m�Fہ����F��1�N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��h�����%�0�u�&�>�3�������KǻN��*ڊ�`�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h_�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF��G1�����1�m�l�u�?�3�}���Y���F�N��U���u�u�%�e�f���������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����H���G��d��U���u�u�u�u�w�}�W���YӖ��lW��V�����'�2�i�u���B���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��h����Y����T��E�����x�_�u�u���B�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��E��
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m�Fځ�	����O�C��U���u�u�u�u�w�}�W���YӖ��lW��G��U��%�e�d�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����d�4�
�9��/�Ͽ�
����C��R��U���u�u�%�e�f�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR�����ߊu�u�u�u�w�}�W���Y���F��1�����9�
�'�2�k�}�(߁�&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�F����ƭ�@�������{�x�_�u�w��(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m�F���&����O��_�����u�u�u�u�w�}�W���Y����9��R	��Hʥ�e�d�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*؊�%�#�1�%�2�}����Ӗ��P��N����u�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��E���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�m�n�}����s���F�N��U���u�u�u�u�'�m�E���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lV��h�����%�0�u�h�'�m�E���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�g�o����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��G���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�I�ԓ�A��S��*ڊ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����9�
�'�2�6�.��������@H�d��Uʥ�e�f�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�f�|�#�8�W���Y���F�N��U���u�u�u�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����O����[��=N��U���u�u�u�u�w�}�W���Y���� 9��h��*���2�i�u�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�f�'�8�W�������A	��D�X�ߊu�u�
�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h]�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�e�f�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(߁�&����Z�G1��F�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��h�����%�0�u�&�>�3�������KǻN��*ڊ�
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����m�l�u�=�9�W�W���Y���F�N��U���u�%�e�a�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��Y����l�N��U���u�u�u�u�w�}�WϮ�I�ғ�C9��S1�����h�%�e�a�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�'�0�<����Y����V��C�U���%�e�a�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�m�C��������hZ�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����9��h��*���2�4�&�2�w�/����W���F�G1��@���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lS��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�e�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�&����_��E��I���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����`�%�0�u�$�4�Ϯ�����F�=N��U���
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����`�4�
�9�~�t����Y���F�N��U���u�u�u�
������E�Ƽ�9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�I�Г�C9��S1�����&�<�;�%�8�8����T�����hX�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}��������T9��S1�L���=�;�_�u�w�}�W���Y���F�N�����c�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�f�}����s���F�N��U���u�u�u�u�'�m�A���&����C��R�����c�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*܊�'�2�4�&�0�}����
���l�N��E���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&Ź��V�
N��*���&�
�#�c�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*܊�%�#�1�|�w�5��ԜY���F�N��U���u�%�e�c�'�8�W��	�֓�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����N����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*݊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�d�e�w�5��ԜY���F�N��U���u�u�u�%�g�j��������V�
N��E���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h^��*���2�4�&�2�w�/����W���F�G1��B���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(߁�&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h^��*���#�1�|�u�?�3�}���Y���F�N��U���%�e�b�%�2�}�JϮ�I����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(ׁ�	����l��PN�����u�'�6�&�y�p�}���Y����9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������l^��N�����u�u�u�u�w�}�W���Y���F��h^��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�l�u�?�3�}���Y���F�N��U���u�u�%�e�o�<�(���&����Z�G1��M���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����hV�����4�&�2�u�%�>���T���F��1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(ׁ����F��h�����#�c�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������hV�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e�m�%�0�w�`����A���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(�������A��V�����'�6�&�{�z�W�W���&ù��R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�m�N���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��-�������� _�C��U���u�u�u�u�w�}�W���Y�����hW�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����d�m�u�=�9�W�W���Y���F�N��U���u�%�e�l�6��������F��1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��h��ʴ�&�2�u�'�4�.�Y��s���C9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��h�����|�u�=�;�]�}�W���Y���F�N�����l�%�0�u�j�-�G��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
�f�<�(���&������^	�����0�&�u�x�w�}���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�d��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����J����[��=N��U���u�u�u�u�w�}�W���Y����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�D���=�;�_�u�w�}�W���Y���F�N����
�%�#�1�'�8�W��	����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p���&������^	�����0�&�u�x�w�}���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���d�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��F���&����O��_�����u�u�u�u�w�}�W���Y����l��PN�U���d�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h_�����9�
�'�2�6�.��������@H�d��Uʥ�d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��\�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��h��*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�g�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&�ԓ�C9��S1�����h�%�d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�d�
�'�2�6�.��������@H�d��Uʥ�d�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N����
�%�#�1�~�}����s���F�N��U���u�u�%�d��/���Y����l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ށ�	����l��PN�����u�'�6�&�y�p�}���Y����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�l��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lW��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��Uʥ�d�4�
�9��/���Y����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����	����R��P �����&�{�x�_�w�}�(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ۊ�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�f�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����Z�G1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lV��G1�����0�u�&�<�9�-����
���9F���*ڊ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������C9��P1����l�u�=�;�]�}�W���Y���F�N��U���%�`�e�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��N�������9F�N��U���u�u�u�u�w�}�W���&ù��l��h����u�
�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�`�e�%�0�w�.����	����@�CךU���
�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lV��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`�e�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u���(������C9��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�9��h��*���2�4�&�2�w�/����W���F�G1��Dڊ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y���R��^	�����f�|�!�0�w�}�W���Y���F�N��U���u�
�
�e�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��l��A�����u�h�%�`�f��������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`�d��/�Ͽ�
����C��R��U���u�u�%�`�f���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h[��E���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��m���������YNךU���u�u�u�u�w�}�W���&ƹ��l��PN�U���
�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�`�d��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�H����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��Dۊ�%�#�1�%�2�}�JϮ�L����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����H¹��V��D��ʥ�:�0�&�u�z�}�WϮ�L����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�d�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ƹ��l��A��\���=�;�_�u�w�}�W���Y���F�G1��Dۊ�'�2�i�u���F�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�e�<�(���&������^	�����0�&�u�x�w�}����H����l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�l�(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u�6���������
O��_�����u�u�u�u�w�}�W���Y���C9��\�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����g�m�u�=�9�W�W���Y���F�N��U���u�%�`�d��-����	����[��h[��G���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h_�����u�&�<�;�'�2����Y��ƹF��h[��G���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�K����TF������!�9�d�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��D؊�%�#�1�|�w�5��ԜY���F�N��U���u�%�`�d��/���Y����T��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&�Փ�C9��S1�����&�<�;�%�8�8����T�����h_�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ӓ� 9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Yۇ��@��U
��M��u�=�;�_�w�}�W���Y���F�N��Uʥ�`�d�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�@������F�N��U���u�u�u�u�w�}����H����l��h����u�
�
�f�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�f�%�2�}����Ӗ��P��N����u�
�
�f�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��]�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`�d��-����P�Ƹ�V�N��U���u�u�u�u�w�}����H����V�
N��@��n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�*���#�1�%�0�w�.����	����@�CךU���
�
�a�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�m�n�}����s���F�N��U���u�u�u�u�'�h�Fہ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������P�C��U���u�u�u�u�w�}�W���Y�����h_�����9�
�'�2�k�}�(ځ�M����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���	����R��P �����&�{�x�_�w�}�(ځ�M����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`�d�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����Hǹ��l��G�����u�u�u�u�w�}�W���Y�����h_�����u�h�%�`�f�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�`�d�
�'�+�����ƭ�@�������{�x�_�u�w��(�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�b�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�%�$�:����A���G��d��U���u�u�u�u�w�}�W���YӖ��lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�`�4��1�(������C9��[�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��h��ʴ�&�2�u�'�4�.�Y��s���C9��[�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�h�Fځ����F��h�����#�c�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����9�|�|�!�2�}�W���Y���F�N��U���
�
�`�%�2�}�JϮ�L����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�B�������W9��R	�����;�%�:�0�$�}�Z���YӖ��lW��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��D���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�l�|�#�8�W���Y���F�N��U���u�u�u�
����������TF���*ۊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����u�&�<�;�'�2����Y��ƹF��h[��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�B���	����[��G1�����9�d�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�'�0�a�W���&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h�E���&����C�������%�:�0�&�w�p�W���	�ӓ�l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(݁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�<�(���&����U�����ߊu�u�u�u�w�}�W���Y���F��1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�e�|�!�2�}�W���Y���F�N��U���u�u�
�
��-����	����[��h[��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��1�����&�<�;�%�8�8����T�����h\�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�h�E��������T�����d�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�'�2�k�}�(ځ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�b�n��������V��D��ʥ�:�0�&�u�z�}�WϮ�L�Փ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u�6���������
O��_�����u�u�u�u�w�}�W���Y���C9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����d�|�!�0�w�}�W���Y���F�N��U���u�
�
�
�'�+���������h]�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��G��U���<�;�%�:�2�.�W��Y����lS��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�n����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��V�����|�!�0�u�w�}�W���Y���F�N��*ߊ�
�'�2�i�w��(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`�c�<�(���&������^	�����0�&�u�x�w�}����M����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����lS��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����9��R	�����;�%�:�0�$�}�Z���YӖ��lR��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�`�c�-����DӇ��P	��C1��D܊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����9��h��\���!�0�u�u�w�}�W���Y���F���*ފ�'�2�i�u���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`�`�6���������@��YN�����&�u�x�u�w�-�B�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����J����[��=N��U���u�u�u�u�w�}�W���Y����9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��F���!�0�u�u�w�}�W���Y���F�N��U���
�
�%�#�3�-����DӖ��lS��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ��C�������%�:�0�&�w�p�W���	�ӓ�l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�`�`�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ƹ��R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h[��*���2�i�u�
��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�`�c�4��1�(���Ӈ��Z��G�����u�x�u�u�'�h�A���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ƹ��R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ߊ�
�%�#�1�'�8�W��	�ӓ�l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&Ź��V��D��ʥ�:�0�&�u�z�}�WϮ�L�Г�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�`�c�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&Ź��l��G�����u�u�u�u�w�}�W���Y�����hX�����i�u�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�`�b�4�
�;���������]F��X�����x�u�u�%�b�j��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����4�
�<�
�3��D�������9F�N��U���u�u�u�u�w�}�W���&Ĺ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��]�����u�u�u�u�w�}�W���Y���F���*݊�%�#�1�%�2�}�JϮ�L�ѓ�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ځ�&������^	�����0�&�u�x�w�}����N����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`�b�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�&����_�N�����u�u�u�u�w�}�W���Y����lS��h����u�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����m�4�
�9��/�Ͽ�
����C��R��U���u�u�%�`�o�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ځ�&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lT��N�����u�u�u�u�w�}�W���Y���F��h[��*���#�1�%�0�w�`����A����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(ׁ�����@��YN�����&�u�x�u�w�-�B���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����m�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(ׁ�	����O�C��U���u�u�u�u�w�}�W���YӖ��l^��E��I���
�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��@���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�`�l�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^�����<�
�1�
�d�t����Y���F�N��U���u�u�u�u�w��(ց�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������W�C��U���u�u�u�u�w�}�W���Y�����hW�����1�%�0�u�j�-�B�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(���Ӈ��Z��G�����u�x�u�u�'�h�N�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��@���%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���(������F��R ��U���u�u�u�u�w�}�W���	�ӓ�l��PN�U���
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��E���
�9�
�'�0�<����Y����V��C�U���%�b�e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*ڊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F��*���
�1�
�f�~�)����Y���F�N��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��h�����%�0�u�h�'�j�G���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�`�m����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��E���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�N�֓�A��S��*݊�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�*���#�1�%�0�w�.����	����@�CךU���
�
�e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�m�n�}����s���F�N��U���u�u�u�u�'�j�F߁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������R�C��U���u�u�u�u�w�}�W���Y�����h_�����9�
�'�2�k�}�(؁�I����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���	����R��P �����&�{�x�_�w�}�(؁�I����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b�d�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����Hù��l��G�����u�u�u�u�w�}�W���Y�����h_�����u�h�%�b�f�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b�d�
�'�+�����ƭ�@�������{�x�_�u�w��(�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�f�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�%�$�:����A���G��d��U���u�u�u�u�w�}�W���YӖ��lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�d�4��1�(������C9��_�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��h��ʴ�&�2�u�'�4�.�Y��s���C9��_�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�Fށ����F��h�����#�c�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����9�|�|�!�2�}�W���Y���F�N��U���
�
�d�%�2�}�JϮ�N����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@��&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&�ԓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����	����l��hV�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�g�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�c�t����Y���F�N��U���u�u�u�u�w��(�������W9��R	��Hʥ�b�d�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����d�
�'�2�6�.��������@H�d��Uʥ�b�d�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lW��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�g�4��1�^�������9F�N��U���u�u�u�u�w��(���	����[��hY��G�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��1��*���
�'�2�4�$�:�W�������K��N�����d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1�*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�f�|�#�8�W���Y���F�N��U���u�u�u�
��n��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��h�����%�0�u�h�'�j�F܁�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`�l�(���Ӈ��Z��G�����u�x�u�u�'�j�F܁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�f�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�9��h����u�
�
�f�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�a�4�
�;���������]F��X�����x�u�u�%�`�l�(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�b�d�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�E���=�;�_�u�w�}�W���Y���F�N�����d�
�%�#�3�-����DӖ��lW��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�9��R	�����;�%�:�0�$�}�Z���YӖ��lW��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��i����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��h�����|�u�=�;�]�}�W���Y���F�N�����d�
�'�2�k�}�(؁�M���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���B���&����C�������%�:�0�&�w�p�W���	�ѓ�9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@��&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��Dߊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�a�l�w�5��ԜY���F�N��U���u�u�u�%�`�l�(�������A��S��*݊�`�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���%�0�u�&�>�3�������KǻN��*݊�`�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����d�
�%�#�3�t�W������F�N��U���u�u�u�%�`�l�(������C9��[�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����9��h��*���2�4�&�2�w�/����W���F�G1��D���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lW��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�D������F�N��U���u�u�u�u�w�}����H����E
��G��U��%�b�d�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�'�2�6�.��������@H�d��Uʥ�b�d�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�W������F�N��U���u�u�u�%�`�l����Y����lQ��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��R��[
�����4�&�2�u�%�>���T���F�� 1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Q����Z��S
��F���!�0�u�u�w�}�W���Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�d�o�W������F�N��U���u�u�u�u�w�-�@�������W9��R	��Hʥ�b�g�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�
�'�2�4�$�:�W�������K��N�����g�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*݊�
�%�#�1�~�}����s���F�N��U���u�u�%�b�e�-����DӖ��lT��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����l��h��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N�Փ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����	����l��hV�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�f�f�}����s���F�N��U���u�u�u�u�'�j�D���&����C��R�����f�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*ي�'�2�4�&�0�}����
���l�N��B���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����V�
N��*���&�
�#�c�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*ي�%�#�1�|�w�5��ԜY���F�N��U���u�%�b�f�'�8�W��	�ѓ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(؁�&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����M����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*ފ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�f�e�w�5��ԜY���F�N��U���u�u�u�%�`�i��������V�
N��B���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hY��*���2�4�&�2�w�/����W���F�G1��A���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*���#�1�|�u�?�3�}���Y���F�N��U���%�b�a�%�2�}�JϮ�N����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(ځ�	����l��PN�����u�'�6�&�y�p�}���Y����9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������l^��N�����u�u�u�u�w�}�W���Y���F��hY��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�f�l�u�?�3�}���Y���F�N��U���u�u�%�b�b�<�(���&����Z�G1��@���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h[�����4�&�2�u�%�>���T���F�� 1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(ځ����F��h�����#�c�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h[�����1�|�u�=�9�W�W���Y���F�N��Uʥ�b�`�%�0�w�`����L���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(�������A��V�����'�6�&�{�z�W�W���&Ĺ��R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�A���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��-�������� _�C��U���u�u�u�u�w�}�W���Y�����hX�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����f�m�u�=�9�W�W���Y���F�N��U���u�%�b�c�6��������F�� 1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��h��ʴ�&�2�u�'�4�.�Y��s���C9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��h�����|�u�=�;�]�}�W���Y���F�N�����c�%�0�u�j�-�@��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������TF��D��U���6�&�{�x�]�}�W���&Ĺ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�j��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����b�u�=�;�]�}�W���Y���F�N��U���%�b�b�4��1�(������C9�� 1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lQ��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��lQ��G1�����u�=�;�_�w�}�W���Y���F�N��B���%�0�u�h�'�j�@�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��-����	����R��P �����&�{�x�_�w�}�(؁�&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b�o�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�%�$�:����A���G��d��U���u�u�u�u�w�}�W���YӖ��l^��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��A��u�=�;�_�w�}�W���Y���F�N��Uʥ�b�m�4�
�;�����E�Ƽ�9��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�l��PN�����u�'�6�&�y�p�}���Y����9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
��/���Y����\��h��C��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ѓ�l��A��\���=�;�_�u�w�}�W���Y���F�G1��M���0�u�h�%�`�e�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(ց�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b�l�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�%�&�0�?���@�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�@���=�;�_�u�w�}�W���Y���F�N�����l�4�
�9��/���Y����
9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�N�ߓ�A��V�����'�6�&�{�z�W�W���&Ĺ��C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�
�%�:�K���	����@��A_��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N�ߓ�C9��SG��U���;�_�u�u�w�}�W���Y���F�� 1�����u�h�%�b�n�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�%�#�3�-����
������T��[���_�u�u�
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�m�n�}����s���F�N��U���u�u�u�u�'�d��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�
9��h��*���2�i�u�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�l�%�0�w�.����	����@�CךU���
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ߓ�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��L���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�'�0�a�W���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�<��4�1���5����@9��P1�Fʴ�&�2�u�'�4�.�Y��s���Z*��^1�����:�
�
�0��d�(�������A	��N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�<�u�4��4�(���&����F��R ��U���u�u�u�u�w�}�W�������l ��h"�����'�2�c�f�k�}�;���&����	��h_�����d�e�%�n�w�}�W���Y���F��[��U´�
�<�
�1��l�^Ϫ���ƹF�N��U���u�u�u�u��1�(���&����l��R	��L���h�4�
�:�$��ځ�B���F�N��U���u�;�u�3�]�}�W���Y���V��^����u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����;�u�:�}�'�.��������O�C�����u�u�u�u�w�}�W���&����r��B��L���'�2�g�f�w�`��������A��C1�*ڊ� �l�e�%�l�}�W���Y���F���*���9�'��!�c��G������� F���*���9�'��!�c�����/����S��G]��Eʱ�"�!�u�e�l�}�W���Y���F���*���9�'��!�c��F�������F���*���9�'��!�c�����/����S��G]��Dʱ�"�!�u�d�l�}�W���Y���F���*���9�'��!�c��E������� F���*���9�'��!�c�����/����S��G]��Gʱ�"�!�u�g�l�}�W���Y���F���*���9�'��!�c��D�������F���*���9�'��!�c�����/����S��G]��Fʱ�"�!�u�f�l�}�W���Y���F���*���9�'��!�c��C������� F���*���9�'��!�c�����/����S��G]��Aʱ�"�!�u�a�l�}�W���Y���F���*���9�'��!�c��B�������F���*���9�'��!�c�����/����S��G]��@ʱ�"�!�u�`�l�}�W���Y���F���*���9�'��!�c��(���&����Z�V������'� �
�n�)����&����^��F����!�u�|�_�w�}�W���Y���F��E1�����'� �
�l�e�/���M�����h������!�a�
�2�-�!���&����CU�
�����g�n�u�u�w�}�W���Y����A��X�����!�a�
�
�2��E��E�ƭ�A9��X�����
�l�!�8�����A���� F��@ ��U���_�u�u�u�w�}�W���Y����Q	��v�� ���l�a�'�2�e�h�W������\	��E����
�0�%��1��Bׁ�J����\��XN�N���u�u�u�u�w�}�WϿ�����_'��x��Aӊ�
�0�
�g�o�a�W���&����r��B��L���8�
�
� �o�e����Y����G	�UךU���u�u�u�u�w�}��������A)��hZ��C���2�g�c�u�j�<��������|��W������3�
�`��n�AϺ�����O��N��U���u�u�u�u�6�/����8����G9��hY�����g�m�i�u�%���������lR��C��*��� �m�m�%��}�������9F�N��U���u�u�u�'��2����6����
9��E��G��u�h�4�'�5�2�6�������l��G1�����`�
�f�m�3�*����P���F�N��U���u�4�'�7�8�����&�ߓ�l��h\�M��u�'�
�:�;�/�8���Mʹ��^��h��M���%�}�u�:�9�2�N��Y���F�N��U���'�
�:�9�%����&ù��T9��]��Hʴ�'�7�:��%�(�(���I����P��G_�U���u�u�u�u�w�}��������A��C1�*���'�2�g�e�w�`����<����|��W�� ��e�%�}�e�3�*����I��ƹF�N��U���u�u�'�
�8�1��������W��R	��G��i�u�����8���Lʹ��l^��h�D���:�;�:�d�~�W�W���Y���F�N�����:��'� ��l�F݁�����U�
N��*����� �
�n�;�(��&���F��@ ��U��n�u�u�u�w�}�W���YӇ��l��[/��:���`�
�f�'�0�o�F���Dӓ��`#��t:�����
� �m�e�'�u�DϺ�����U�=N��U���u�u�u�u�w�/�(�������F��1�*���
�g�f�i�w�
�$���:����lS��Q��@ڊ�f�d�u�:�9�2�F���s���F�N��U���4�'�7�:��/����H����A��\�U�� �
����(�(�������9��_����!�u�`�n�w�}�W���Y���F��E�����'��!�`������H���F��h=��0��� �
�l�3��h�(��Hӂ��]��G�U���u�u�u�u�w�}��������A��C1�*؊�0�
�d�f�k�}� ���5����F��1��*���
�f�g�1� �)�W���s���F�N��U���4�'�7�:��/����H�Փ�V��X�I��������)�Bց�����l��N�����u�|�_�u�w�}�W���Y���R��U��4��� �
�d�a�%�:�E��Y����d9��{+��:���`�
� �m�g�-�_�������R�=N��U���u�u�u�u�w�/�(�������F��1�����g�b�u�h�"��2���-����_��B1�E���}�u�:�;�8�h�L���Y���F�N��U���
�:�9�'��)�Bށ�&����W��R�� ������ ��d����Lù��P��X����n�u�u�u�w�}�W���YӇ��l��[/��:���`�
�
�0��l�O��Y����v*��c!��*���3�
�`�
�d�j��������l�N��U���u�u�u�4�%�?��������W��h��*��f�i�u����4�������U��^��F��1�"�!�u�~�W�W���Y���F�N�����:��'� ��l�N�������F���&�����!�`��(�O���	����W	��C��\�ߊu�u�u�u�w�}�W�������\
��E!��*���e�'�2�g�`�}�JϿ�����_'��x��@ي�
� �b�a�'�f�W���Y���F�N�����:�9�'��#�h�(�������T��S��*ۊ�;�&�2�d�w�2����H����F�N��U���u�u�4�'�5�2�6�������lW��E��G��u�h�%�d�>�����Hӂ��]��_����u�u�u�u�w�}�W���&����r��B��F��
�0�
�d�d�a�W���&����Z�N�����u�g�n�u�w�}�W���Y�����h������!�`�
�d�/���J�����h�����d�u�:�;�8�l�^�ԜY���F�N��Uʴ�'�7�:��%�(�(���Hǹ��T9��]��Hʥ�d�<�
�<��i��������]ǻN��U���u�u�u�u�%���������lS��[�����d�m�i�u����������W	��C��@��u�u�u�u�w�}�W�������\	��E�����
�
�0�
�g�e�K���&¹��l��_�����:�d�n�u�w�}�W���Y�����h������!�`�
��8�(��J���C9��^ �����u�:�;�:�e�f�W���Y���F�N�����:�9�'��#�h�(܁�����^�
N��D���
�<�}�u�8�3���B���F�N��U���u�'�
�:�;�/�8���L����A��^�U��%�d�<�
�>�u�W������]ǻN��U���u�u�u�u�%���������lS��1����l�u�h�%�f�4�(���Q�ƨ�D��[����u�u�u�u�w�}�W���&����r��B��F���'�2�g�e�w�`��������TN��S�����|�_�u�u�w�}�W���Y�ƭ�A9��X�����
�f�b�'�0�o�G���DӖ��l��D��Bʱ�"�!�u�|�]�}�W���Y���F�V������'� �
�d�e����K����[��h_�����2�m�1�"�#�}�^�ԜY���F�N��Uʴ�'�7�:��%�(�(���@����lT��N�U���
�;�&�2�n�9� ���Y����F�N��U���u�u�7�:���3���2����F��1�I���
�g�'�4��8����&����CT��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D��ۊ�u�u�-�!�8�9�(���H����CT�V ��]���
� �d�g��l�JϿ�&����G9��1��\���=�;�u�u�w�}�W���Y����A��C1�����:�
�b�d��m����N�����h��3����:�
�b�g�;�(��O����9F�N��U���u�u�u�'��)�1���5����_��1�*���f�c�i�u�%���������C9��h^�� ��l�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h_�����}�%�6�;�#�1�F��DӃ��G��SY�� ��d�
�g�u�9�}��������P��N�����:�&�
�#��t�^Ϫ����F�N��U���u�4�'�9��2�(���	����S��1��*��u�h�4�'�;���������9��Q��G���%�n�u�u�w�}�W���Y����A��C1�����:�
�l�d��l����M�����h��3����:�
�l�g�;�(��K����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������]��[��E��0�<�6�;�`�;�(��M������F�����
�d�c�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����_��X�����g�
�`�d��(�E��E�ƭ�A9��h(��*���%�g�
�
�"�l�Oف�K���F�N��U���u�4�'�9��2�(���	����S��1��*��u�h�4�'�;���������
9��Q��G���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U´�
�:�&�
�!��W�������]��Q��D���%�|�4�1��0�(���H����CW������!�9�a��~�}����Y���F�N��U���'�
�!��%�����N����U��B1�A��u�'�
�!��/�;���&�ѓ�l ��\�*��_�u�u�u�w�}�W���Y����_��X�����g�
�`�d��(�D��E�ƭ�A9��h(��*���%�g�
�
�"�l�N݁�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��h^��U���!�:�1�
�"�l�Fہ�K�ƭ�WF��Z�� ��g�
�d�h�6�����&����vO������u�u�u�u�w�}�WϿ�����u	��{��*���d�
�a�3��e�W������G9��E1�����b�e�3�
�e�k���Y���F�N��U���'�
�!��%�����@����R��B1�G��u�'�
�!��/�;���&�ߓ�l ��\�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�d�g�`��������l ��_�*��u�;�u�:��)����&����l��
N��*���&�
�#�
�~�}��������^��B1�G܊�d�h�4�
�8�.�(���&���R��Y��]���
� �d�g��l�JϿ�&����G9��1��\ʴ�1�;�!�}�:����KŹ��[��G1�����9�a��|�6�9����Q����U��\�����u�%�6�;�#�1�C���PӇ����F�����
�d�c�%�w�}��������ER��G�����:�}�!�%�1��F���	���R��X ��*���
�|�u�;�w�2�_Ǫ�	����W��h�Hʴ�
�:�&�
�!��^����Ƣ�GN��Z�� ��g�
�d�h�6�����&����O�V �����}�8�
� �f�o�(��DӇ��P	��C1��A���|�4�1�;�#�u��������9��S�����;�!�9�a�c�t�������G��Q��D���%�u�u�%�4�3����M����� ��]¡�%�3�
�d�a�-�W���	����@��AZ��\���;�u�:�}�#�-����H�Г�F�V�����
�#�
�|�w�3�W���Qے��l ��_�*��h�4�
�:�$��ہ�P���G��=N��U���u�u�u�u�w�/�(���?����\	��Y��@��
� �g�g�k�}��������l*��G1�*ڊ� �d�m�
�e�W�W���Y���F�N�����
�:�
�:�'�o�(���Hƹ��lU��R�����9�
�:�
�8�-�Eց�&����_��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����#�
�u�u�/�)����&����W��G\�����}�8�
� �f�o�(��DӇ��P	��C1��A��|�u�=�;�w�}�W���Y���F��E�����'��:�
�`�l�(ށ�����Z�V�����:�
�:�%�e��(���H����CT��N��U���u�u�u�u�6�/��������\��1�*ۊ� �f�e�i�w�/�(���?����\	��W��*���d�l�
�g�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʴ�1�}�%�6�9�)����I����K��X ��*���d�d�
�g�w�3�WǪ�	����W��h�Hʴ�
�:�&�
�!��^�������F�N��U���u�u�4�'�;���������9��h\�� ��e�i�u�'��)�1���5����Q��h��D��
�g�_�u�w�}�W���Y���R��[�����:�%�g�
�b�o����I�����h��3����:�
�l�g�;�(��K����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������]��[��E��0�<�6�;�`�;�(��M������F�����
�d�c�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����_��X�����g�
�`�f�1��C���DӇ��l
��q��9���
�b�e�3��o�A���B���F�N��U���u�'�
�!��/�;���&�ߓ�9��Q��E���h�4�'�9��2�(���	����9��h_�G���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�#��}�W�������9��h_�A���|�4�1�}�:����KŹ��[��G1�����9�a�a�|�w�5����Y���F�N��U���
�!��'��2�(���Hƹ��U��V��Hʴ�'�9�
�:��2���&ù��lW��1��N���u�u�u�u�w�}�WϿ�����u	��{��*���d�
�
� �d�o�K�������l ��h"����
�
� �d�n��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������lV������1�
� �d�f��E�������^��B1�G܊�d�h�4�
�8�.�(���&�����Yd��U���u�u�u�u�w�<����&����	��h\��Dߊ�
� �g�g�k�}��������l*��G1�*ڊ� �d�m�
�e�W�W���Y���F�N�����
�:�
�:�'�o�(���L���� W��S�����!��'��8��N�������
T��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�;���Y������T�����d�e�h�0�>�>��������R��G�����!�%�3�
�f�k����Y����\��h��*���|�!�0�_�w�}�W���Y���F��E1��*���
�:�%�g��h�A���&����[��E�����'��:�
�`�m����K�Г�]ǻN��U���u�u�u�u�%���������C9��h_��C���
�g�u�h�6�/��������\��1�����g�g�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$��ށ�Y�Ʃ�Z��Y
�����d�a�%�|�6�9�_���&����T��G_��U���6�;�!�9�c�j�^�����ƹF�N��U���u�u�'�
�#���������lW�� 1��*��u�h�4�'�;���������9��Q��G���%�n�u�u�w�}�W���Y����A��C1�����:�
�l�d�����M���R��[�����:�%�g�
��(�F��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��A_��U���-�!�:�1��(�F��&���R����*���d�g�
�d�j�<�(���
����9��G�����u�u�u�u�w�}�W�������G9��E1�����b�d�
�
�"�o�C��Y����_��X�����g�
�
� �f�e�(��s���F�N��U���4�'�9�
�8�����Kʹ��l^��B1�M��u�'�
�!��/�;���&�ߓ�l ��\�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�d�g�`��������l ��_�*��u�;�u�!�'�;�(��O����F��h�����#�
�|�|�#�8�}���Y���F�N�����9�
�:�
�8�-�E؁�L�ߓ�F9��N�U���
�!��'��2�(���I����T��h����u�u�u�u�w�}�W���&����\��X��Gӊ�`�l�3�
�d�}�JϿ�����u	��{��*���e�3�
�g�e�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�u�;�u�6�����&����F�R�����b�3�
�d�c�-�^Ͽ��θ�C9��h_�C���u�u�%�6�9�)����I���G��=N��U���u�u�u�u�w�/�(���?����\	��Y��@���
�f�u�h�6�/��������\�� 1�����g�c�%�n�w�}�W���Y���F��E�����'��:�
�n�l�(���K���F��E1��*���
�:�%�g�����@����l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӒ����CN�����}�%��
�$�t�����ƿ�R��Z�����u�x�u�u�6��$�������Z��G��U���'�6�&�u�6��$����ƭ�l�������7�1�c�a�w�%����Ĺ��lW��1��\���u�7�2�;�w�}�W�������R��d1��ʼ�_�u�u�u�w�}�W���Ӈ��`2��C_�����u�k�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X�����2�7�1�c�c�t�W������F�N��U���u�u�u�%������DӇ��`2��C\�����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=�����3�8�e�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��Q��D��u�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	�������!�9�d�e�j�8�����ѓ�F9��Z��G���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����l ��h_�U���u�u�u�u�w�}������ƹF�N��U���=�;�:�=�%�}�I���Y���F�N��U���%��
�&�w�`�U���B���F���U���0�_�u�u�9�}����
��ƓF�C�����;�u�&�<�9�-����
���9F������
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������F��^�����3�
�d�a�'�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Y������T�����d�e�h�0�>�>��������R��G��\ʡ�0�u�u�u�w�}�W�������]�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�3�3�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�����ƭ�@�������{�x�_�u�w�-����&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�]�}�W������F�N��U���:�}�4�
�8�.�(�������F��h�����u�;�u�4��2��������F�V�����&�$��
�#�����P����[��=N��U���u�u�u�%�>�1�W������]��[����_�u�u�u�w�1��ԜY���F�N��*���0�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�0�1�w�.����	����@�CךU���%�'�4�,�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���!�:�1�
�"�l�Fہ�K���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����:�&�
�#��}�W�������9��h_�A���|�|�u�=�9�W�W���Y���F��h�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W�������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����e�4�&�2�w�/����W���F�V�����1�
�e�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�e�`�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��W�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��M���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�N��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l_��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�d�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�@Ͽ�
����C��R��U���u�u�4�
�>�����KĹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(߁�I����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����V��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�f�w�.����	����@�CךU���%�&�2�7�3�l�A���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�g�l�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��]�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����H¹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����d�`�4�&�0�}����
���l�N��*���
�1�
�a��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�g�6�����Y����V��=N��U���u�u�u�u�w�-��������S�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���E���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��A��4�&�2�u�%�>���T���F��h��*���
�a�a�4�$�:�(�������A	��D�����2�6�0�
��.�E������V��T��B���
�d�a�%�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���O���N��G1�����9�2�6�d�j�<�(���&����l5��D�����d�u�;�u�6�����&����F�R�����b�3�
�d�c�-�^��Y����]��E����_�u�u�x�w�-��������R��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��[�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��]�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�b�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��E��
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����O�ƭ�@�������{�x�_�u�w�-��������U��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�f�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�EϿ�
����C��R��U���u�u�4�
�>�����N����@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(߁�L����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����S��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�m�6�.��������@H�d��Uʴ�
�<�
�1��e��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����H���N��h-�����e�1�"�!�w�t�JϿ�&����G9��1�N���u�0�1�%�8�8��Զs���K��G1�����1�d�d�4�$�:�W�������K��N�����<�
�1�
�o���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�f�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��^�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��E���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�G��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��lW��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�l�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�OϿ�
����C��R��U���u�u�4�
�>�����I˹��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ځ�&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��G��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ӓ�l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�d�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�j��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�`�d�<�(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(܁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��G��4�&�2�u�%�>���T���F��h��*���
�g�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����K���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`�a�6�����B����������n�_�u�u�z�}��������lT�������%�:�0�&�w�p�W�������T9��S1�@���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�e�h�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ߊ�
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������R��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ӓ�l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�a�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�e�n�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(؁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�F��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�L�ѓ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�c�u�&�>�3�������KǻN�����2�7�1�g�e�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�`�m�6�����Y����V��=N��U���u�u�u�u�w�-��������T�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Dʴ�&�2�u�'�4�.�Y��s���R��^	�����b�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ߊ�
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`�l�4��1�^��Y����]��E����_�u�u�x�w�-��������V��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��V�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��^�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�o�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��@��
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����A�ƭ�@�������{�x�_�u�w�-��������_��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ӓ�9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�g�l�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�OϿ�
����C��R��U���u�u�4�
�>�����@˹��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ځ�K����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����T��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�e�w�.����	����@�CךU���%�&�2�7�3�n�@���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�b�l�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��^�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����H����l��G�U���0�1�%�:�2�.�}�ԜY�����D�����f�c�4�&�0�}����
���l�N��*���
�1�
�d��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�a�6�����Y����V��=N��U���u�u�u�u�w�-��������P�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���C���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��G���&�<�;�%�8�8����T�����D�����f�`�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^����d�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����K���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`�d��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Fފ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��hY��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��n�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����e�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� R��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�f�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��h�W�������A	��D�X�ߊu�u�%�&�0�?���K����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��@���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�f�d�4�$�:�W�������K��N�����<�
�1�
�a���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&���� P��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�D���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��Bʴ�&�2�u�'�4�.�Y��s���R��^	�����b�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��E���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�D���D����C9��Y�����6�d�h�%�g�m��������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��V�����u�u�7�2�9�}�W���Y���F������7�1�f�e�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��@���
������T��[���_�u�u�%�$�:����J�ߓ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����L����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����9��h��\��u�u�0�1�'�2����s���F������7�1�f�m�6�.��������@H�d��Uʴ�
�<�
�1��e�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
���������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�b�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b�b�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����J���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��E܊�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��hY��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��m�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����m�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����M����@��YN�����&�u�x�u�w�<�(���&����W��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����
9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�a�`�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������hW�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��o�W�������A	��D�X�ߊu�u�%�&�0�?���M����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��A��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ѓ�9��h��\��u�u�0�1�'�2����s���F������7�1�a�f�6�.��������@H�d��Uʴ�
�<�
�1��n�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��l������ƹF��R	�����u�u�u�u�w�}�W���
����W��]��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�H����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����a�u�&�<�9�-����
���9F������7�1�a�g�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�b�d�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`�l�(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Dʴ�&�2�u�'�4�.�Y��s���R��^	�����`�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*݊�f�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���H�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�f�6�����B����������n�_�u�u�z�}��������lR��V�����'�6�&�{�z�W�W���	����l��hZ�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�w�`�_���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��D���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&�ғ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����c�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�a�}����Ӗ��P��N����u�%�&�2�5�9�C�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�j�Fځ�	����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�a�e�4�$�:�W�������K��N�����<�
�1�
�o���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�n�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��_�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��d�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N����
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����I�ƭ�@�������{�x�_�u�w�-��������V��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	����R��[
��U���7�2�;�u�w�}�W���Y�����D�����`�e�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lW��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�`�w�.����	����@�CךU���%�&�2�7�3�h�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
���������F��P��U���u�u�u�u�w�}��������W9��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(݁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��C��4�&�2�u�%�>���T���F��h��*���
�d�
�&�>�3����Y�Ƽ�\��DF��*���'�y�%�e�g�<�(���&����Z�G1��D���
�9�
�;�$�:�W���&����l��h�����u�
�
�
�'�+����&������hZ�����1�<�
�<�{�-�G�������W9��h��Yʥ�e�c�4�
�;������Ƽ�9��V�����;�&�2�u���(�������]9��PB��*ڊ�
�%�#�1�>����	�֓�9��h��*���&�2�u�
��l��������l��N��E��
�%�#�1�>����	�֓� 9��h��*���&�2�u�
��i��������l��N��E��
�%�#�1�>����	�ד�C9��S1��*���y�%�`�e�6���������F��1�����9�
�;�&�0�}�(ځ�&����_��Y1�����
�
�
�%�!�9��������lS��h�����<�
�<�y�'�h�B���&����Z��^	����c�4�
�9��3����Y����9��h��*���&�2�u�
����������@����*ӊ�%�#�1�<��4�[Ϯ�L����R��[
�����2�u�
�
�f�<�(���&����Z�G1��D؊�%�#�1�<��4�[Ϯ�L����R��[
�����2�u�
�
�c�<�(���&����Z�G1��Dߊ�%�#�1�<��4�[Ϯ�N�֓�C9��S1��*���y�%�b�d�6���������F�� 1�����9�
�;�&�0�}�(؁�&����_��Y1�����
�
�
�%�!�9��������lQ��h�����<�
�<�y�'�j�A���&����Z��^	����b�4�
�9��3����Y����9��h��*���&�2�u�
����������@����*���4�
�9�
�9�.����&Ĺ��l��A�����<�y�%�b�f���������@����*���4�
�9�
�9�.����&Ĺ��l��A�����<�y�%�b�f���������@����*���#�1�<�
�>�q���&����_��Y1�����
�g�4�
�;��������F��P��U���u�u�u�u�w�}��������W9��N�U���
�g�4�
�;���������C9��Y�����6�e�u�'���F���&����Z��^	��U���6�;�!�9�0�>�G����μ�
9��h��*���&�2�h�4��2��������O��EN��*ۊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`�g�<�(���&����Z������!�9�2�6�g�}����&ƹ��R��[
�����2�h�4�
�8�.�(�������	����*؊�%�#�1�<��4�W���	����@��X	��*���:�u�%�`�d�<�(���&����Z������!�9�2�6�g�}����&ƹ��R��[
�����2�h�4�
�8�.�(�������	����*ߊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`�a�<�(���&����Z������!�9�2�6�g�}����&ƹ��R��[
�����2�h�4�
�8�.�(�������	����*Ҋ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`�n�<�(���&����Z������!�9�2�6�g�}����&ƹ��l��A�����<�u�u�%�4�3��������F��F��@��
�%�#�1�>�����Y����\��h�����|�:�u�%�b�l�(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��lW��V�����;�&�2�h�6�����&����P9����]���
�a�4�
�;���������C9��Y�����6�e�u�'���(�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�@�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�@�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�@�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�e�4��1�(���
�����T�����2�6�e�u�%�u�(؁�H����E
��^ �����u�%�6�;�#�1����I�ƣ�N�� 1�*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b�d��-��������TF�V�����
�:�<�
�~�2�WǮ�N����R��[
�����2�h�4�
�8�.�(�������	����*���4�
�9�
�9�.�������]��[����u�'�}�
����������@��
N��*���&�
�:�<��t����	�֓�l��A�����<�u�u�%�4�3��������F��F��E���4�
�9�
�9�.�������]��[����u�'�}�
����������@��
N��*���&�
�:�<��t����	�֓�l��A�����<�u�u�%�4�3��������F��F��E���4�
�9�
�9�.�������]��[����u�'�}�
����������@��
N��*���&�
�:�<��t����	�֓�l��A�����<�u�u�%�4�3��������F��F��E���4�
�9�
�9�.�������]��[����u�'�}�
����������@��
N��*���&�
�:�<��t����	�֓�9��h��*���&�2�h�4��2��������O��EN��*ڊ�d�4�
�9��3����DӇ��P	��C1�����e�u�'�}���E���&����Z��^	��U���6�;�!�9�0�>�G����μ�9��h�����<�
�<�u�w�-��������Z��N��U¥�e�d�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G��&����_��Y1����4�
�:�&��2����PӉ����D����4�
�:�&��2����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Y�����;�%�:�0�$�}�Z���YӇ��@��U
��C���4�&�2�
�%�>�MϮ�������D�����
��&�d�1�0�G���	����l��hX�\���u�7�2�;�w�}�W���Y���F��G1�����1�c�b�i�w�u��������\��h_��U���&�2�6�0��	��������F��SN��´�
�<�
�1��l�^��Y����]��E����_�u�u�x�w�-��������F��D��U���6�&�{�x�]�}�W���
����W��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��V�����u�u�7�2�9�}�W���Y���F������7�1�c�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�j�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(ہ�	����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&ǹ��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����m�c�4�&�0�}����
���l�N��*���
�1�
�d��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Y����G	�G�U���0�1�%�:�2�.�}�ԜY�����D�����m�u�&�<�9�-����
���9F������7�1�m�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Fӊ�&�<�;�%�8�}�W�������R��^	������
�!�
�$��[ϻ�����WQ��B1�Dފ�g�_�u�u�2�4�}���Y���F�N�����<�
�1�
�d�}�J�������]��[����h�4�
�<��.����&����U��G�����:�}�4�
�8�.�(���&���V��T��B���
�d�a�%�~�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����
W��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�d�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ށ�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�m�_�w�}����s���F�^�����<�
�1�
�o�}����s���F�N�����<�
�&�$���ށ�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*ۊ�&�<�;�%�8�}�W�������R��^	�����d�|�u�u�5�:����Y����������7�1�m�c�w�5��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�ƭ�A9��X�����
�l�e�3��d�(��E�ƭ�A9��X�����
�l�!�8�����A����F�N�����u�|�_�u�w�/�(�������F��1�����
� �m�m�'�}�J�ԜY���F��h�����#�c�e�"�2�}����&����|��Y�� ��a�%�}�|�j�z�P������F�N�����<�
�<�n�w�}��������A��C1�*ڊ� �m�c�%�w�`����<����|��W�� ��e�%�}�u�w�}�������9F���*���9�'��!�b��(���N�ғ�F���*���&�2�d�x�f�9� ���Y����F�V�����:�
�:�%�e��(���H����CT�
N�����;�1�
�0�:�n�(���H����CT��Y
�����9�
�:�
�8�-�Eف�����9��G�U���4�'�9�
�8�����Kʹ��U��W�����h�}�:�9�9�9�(�������U��V�����;�u�:�9�;���������9��h_�E���m�n�u�u�5�2�(�������^9��h��D��
�g�i�u�5�2�(��� ���� W��B1�C؊�g�:�u�:�;�1�(���&����lT��Q��D���%�m�n�u�w�?��������V��Y�� ��m�
�g�i�w�?����5����G9��h��D��
�g�:�u�8�1��������\��1��*��m�%�m�n�w�}����&����|��_�� ��c�
�g�i�w�l�W����ο�T�������:�
�:�%�f����Jù��O������<�
�!��%�����A����W��h�\���9�0�w�w�]�}�W�������J)��hX��E���
� �m�m�'�}�J�������v#��v-�� ���!�b�
�u�8�}��������EW��UךU���:�9�-���)�A؁�����l��S��E���
�g�<�
�>�q�������A�=N��U���9�-���#�k�(���A�ғ�F�F������,� �
�`�;�(��&����]��X������!�c�
�#�-����J˹��]ǻN�����-���!�c����O˹��Z�_�����u�&�2�0��
��������\��1��*��e�%�m�u�w�4��������l ��h"����
� �d�b��l�^������D��N�����6�;�b�3��l�C���Y���D��_��]���9�
�:�
�8�-��������[��G1�����9�`�d�|�2�.�W��B�����[�����:�%�d�
�"�l�E߁�K���@��[�����6�:�}�;�>�3�Ƿ�&����\��X�����2�c�f�u�w�3����ۇ��P	��C1��@��|�_�u�u�z�}�(߁�&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�;�&�2�6�.���������T��]���
�
�%�#�3�}�(߁�&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g�m�������G��d��U���u�u�u�%�g�m��������l��R�����e�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
��-��������TF���*ڊ�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h^�����2�4�&�2�w�/����W���F�G1��E���
�<�
�&�>�3����Y�Ƽ�\��DF��E��u�
�
�
�%�:�W���&ù��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��-����PӒ��]FǻN��U���u�u�
�
��3����E�Ƽ�9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��^ �����h�%�e�e�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h^��E���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�e�d��-��������T9��D��*���6�o�%�:�2�.����Hù��l��N��E��
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�*���#�1�|�!�2�}�W���Y���F��h^��E���
�9�
�;�$�:�K���&ù��l��A�����u�u�u�9�2�W�W���Y���F��1�*���#�1�<�
�>�}�JϮ�I����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(߁�I����@��V�����'�6�&�{�z�W�W���&ù��l��D�����2�
�'�6�m�-����
ۖ��lW����*���%�0�y�%�g�l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�e�4�
�;�t�W������F�N��Uʥ�e�d�
�;�$�:�K���&ù��l�N��Uʰ�&�u�u�u�w�}�W���	�֓�9��h��U��%�e�d�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�d�6���������l��^	�����u�u�'�6�$�u�(߁�H����E
����*���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h_�����9�|�u�=�9�W�W���Y���F��1�*���#�1�<�
�>�}�JϮ�I����R��[
�U���u�u�0�&�w�}�W���Y�����h_�����9�
�;�&�0�a�W���&�ד�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�G��&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I����Z��^	�����;�%�:�u�w�/����Q����W�G1��Dۊ�'�2�u�
��l������ƹF��R	�����u�u�u�3��<�(���
����T��N�����d�
�%�#�3�t����Y���F�N��U���
�d�<�
�>�}�JϮ�I����9F�N��U���0�_�u�u�w�}�W���&ù��l��D��I���
�
�d�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h_�����9�
�;�&�0�<����Y����V��C�U���%�e�d�
�'�+����&����R��P �����o�%�:�0�$�-�G��&����_�G1��D؊�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��\�����1�|�!�0�w�}�W���Y�����h_�����9�
�;�&�0�a�W���&�ԓ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��\�����1�<�
�<�w�`����H����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������TF��D��U���6�&�{�x�]�}�W���&�ԓ�]9��P1�����
�'�6�o�'�2����	�֓�J��h^��G���0�y�%�e�f��������F��P��U���u�u�<�u��-��������Z��S��*ڊ�g�4�
�9�~�}����s���F�N�����d�
�;�&�0�a�W���&����F�N�����u�u�u�u�w�}�WϮ�I����Z��^	��Hʥ�e�d�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��]�����1�<�
�<�w�.����	����@�CךU���
�
�f�4��1�(���
����@��Y1�����u�'�6�&���(�������WJ��h^��F���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lV��1��*���|�u�=�;�]�}�W���Y���C9��]�����1�<�
�<�w�`����H����l��d��U���u�0�&�u�w�}�W���Y����lV��1��*���
�;�&�2�k�}�(߁�J����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�F܁�������^	�����0�&�u�x�w�}����H����l��h�����%�:�u�u�%�>����&ù��F��1�*���2�u�
�
�d�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��E��
�%�#�1�~�)����Y���F�N��*ڊ�f�<�
�<�w�`����H��ƹF�N�����_�u�u�u�w�}�W���&�Փ�]9��PN�U���
�f�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lV��1��*���
�;�&�2�6�.��������@H�d��Uʥ�e�d�
�%�!�9��������@��h����%�:�0�&�'�m�Fہ�	����F��1�*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��h�����|�!�0�u�w�}�W���Y����lV��1��*���
�;�&�2�k�}�(߁�M����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��h�����<�
�<�u�j�-�G��&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���C���&����R��P �����&�{�x�_�w�}�(߁�M����@��V�����'�6�o�%�8�8�Ǯ�I������h_�����y�%�e�d��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���4�
�9�|�w�5��ԜY���F�N��E��
�;�&�2�k�}�(߁�M���F�N�����u�u�u�u�w�}����Hǹ��l��R�����d�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�`�4�
�;���������Z��G��U���'�6�&�}���B���&������h_�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lW��V�����u�=�;�_�w�}�W���Y�Ƽ�9��h�����<�
�<�u�j�-�G��&����_��N��U���0�&�u�u�w�}�W���YӖ��lW��V�����;�&�2�i�w��(�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g�l�(���
����@��YN�����&�u�x�u�w�-�G��&����Z��D�����:�u�u�'�4�.�_���&���C9��[�����u�
�
�`�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��Dߊ�%�#�1�|�#�8�W���Y���F���*���<�
�<�u�j�-�G��B���F����ߊu�u�u�u�w�}�(߁�L����@��S��*ڊ�`�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lW��G1�����
�<�u�&�>�3�������KǻN��*ڊ�
�%�#�1�>�����
����l��TN����0�&�%�e�f�<�(���UӖ��lW��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&¹��l��G�����_�u�u�u�w�}�W���&¹��l��h�����i�u�
�
��-����s���F�R��U���u�u�u�u�w�-�G�������W9��h��U��%�e�d�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����d�<�
�<�w�.����	����@�CךU���
�
�
�;�$�:��������\������}�
�
�y�'�m�F�������lV��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G�������WO�C��U���u�u�u�u�w�-�G�������TF���*��u�u�u�u�2�.�W���Y���F���*ۊ�;�&�2�i�w��(ށ�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�e�g�4�
�;�����Ӈ��Z��G�����u�x�u�u�'�m�E���&����Z��^	�����;�%�:�u�w�/����Q����9��h��Yʥ�e�g�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*؊�%�#�1�|�#�8�W���Y���F���*؊�%�#�1�<��4�W��	�֓�l��A�����u�u�u�9�2�W�W���Y���F��1�����9�
�;�&�0�a�W���&����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(݁�������^	�����0�&�u�x�w�}����K����@��V�����'�6�o�%�8�8�Ǯ�I���C9��1�����%�e�g�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����9�|�u�=�9�W�W���Y���F��1�����<�u�h�%�g�o�}���Y���V
��d��U���u�u�u�%�g�o���������h\�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(߁�&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�;�&�2�6�.���������T��]���
�
�%�#�3�}�(߁�&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g�n�������G��d��U���u�u�u�%�g�n��������l��R�����f�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
��-��������TF���*ي�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h]�����2�4�&�2�w�/����W���F�G1��F���
�<�
�&�>�3����Y�Ƽ�\��DF��E��u�
�
�
�%�:�W���&����l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��-����PӒ��]FǻN��U���u�u�
�
��3����E�Ƽ�9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��^ �����h�%�e�f�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h^��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
�'�+����&����R��P �����o�%�:�0�$�-�G�������WJ��h^��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��V�����;�&�2�i�w��(ہ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�֓�l��A�����<�u�h�%�g�i��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�e�a�>�����
������T��[���_�u�u�
����������Z��G��U���'�6�&�}���[Ϯ�I�ғ�A����*ފ�%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�֓�l��A��\ʡ�0�u�u�u�w�}�W���	�֓�l��D��I���
�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�;�$�:�K���&ù��C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e�b�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I�ӓ�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����9�y�%�e�b�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�%�!�9���������h[�����1�_�u�u�w�}����s���F�N�����`�4�
�9��3����E�Ƽ�9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��Z��^	�����;�%�:�0�$�}�Z���YӖ��lS��Y1�����&�2�
�'�4�g��������lV��N��E���%�0�y�%�g�h������ƹF��R	�����u�u�u�3��<�(���
����T��N�����`�4�
�9�~�}����s���F�N�����`�<�
�<�w�`����L���F�N�����u�u�u�u�w�}����L����@��S��*ڊ�
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��h��*���&�2�4�&�0�}����
���l�N��E���4�
�9�
�9�.����
����C��T�����&�}�
�
��-����Y����9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����O����E
��N�����u�u�u�u�w�}����O����E
��^ �����h�%�e�c�6����Y���F��[�����u�u�u�u�w��(ف�	����l��D��I���
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�
�;�&�2�6�.��������@H�d��Uʥ�e�c�<�
�>���������PF��G�����%�e�c�u���(����Ƽ�9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(ف�	����O��_�����u�u�u�u�w��(ف�����Z�G1��C�ߊu�u�u�u�;�8�}���Y���F�G1��C���
�<�u�h�'�m�A�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(�������]9��P1�����
�'�6�o�'�2����	�֓�l��A��U���
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��B���
�9�|�u�?�3�}���Y���F�G1��B���
�9�
�;�$�:�K���&ù��R��[
�U���u�u�0�&�w�}�W���Y�����hY�����1�<�
�<�w�`����N����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�@���&����R��P �����&�{�x�_�w�}�(߁�&����Z��D�����:�u�u�'�4�.�_���&����lV��h�����
�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������hY�����1�|�!�0�w�}�W���Y�����hY�����2�i�u�
��f�W���Y����_��=N��U���u�u�u�
���������C9�� 1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�G�������W9��h��U���<�;�%�:�2�.�W��Y����lV��h�����<�
�<�
�$�4��������C��R�����m�4�
�9�{�-�G�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
����������[��=N��U���u�u�u�
����������@��S��*ڊ�
�%�#�1�]�}�W���Y����l�N��U���u�%�e�m�6���������Z�G1��M���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��1��*���u�&�<�;�'�2����Y��ƹF��h^��*���&�2�4�&�0�����CӖ��P����*���%�e�m�%�2�q����A����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�e�m�6�����Y����l�N��U���u�%�e�m�>�����DӖ��l^��N��U���0�&�u�u�w�}�W���YӖ��l^��Y1����u�
�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�����9�
�;�&�0�<����Y����V��C�U���%�e�l�4��1�(���
����@��Y1�����u�'�6�&���(ց�	����F��1�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l_��G1�����!�0�u�u�w�}�W���YӖ��l_��G1�����
�<�u�h�'�m�N���&����9F�N��U���0�_�u�u�w�}�W���&ù��R��[
�����2�i�u�
����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
�9�.�Ͽ�
����C��R��U���u�u�%�e�n�4�(���&����T��E��Oʥ�:�0�&�%�g�d�W���&ʹ��V�G1��L���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��R��[
��U���;�_�u�u�w�}�W���&ù��Z��^	��Hʥ�e�l�_�u�w�}�W������F�N��Uʥ�e�l�<�
�>�}�JϮ�I�ߓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�e�i�u��8����L����F9��Z��D��_�u�u�x�'�l�(�������@��YN�����&�u�x�u�w�-�F߁�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�3�8�f�}��������U��_�����u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����u�;�u�:��<�(���
����9��
N�����;�b�3�
�f�i����P�Ƹ�V�N��U���u�u�%�d��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���e�4�
�9�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u��l��������l�������%�:�0�&�w�p�W���	����R��[
�����2�4�&�2��/���	����@��h_�����9�y�%�d��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�d�
�%�#�3�t����Y���F�N��U���d�4�
�9��3����E�Ƽ�W��G1���ߊu�u�u�u�;�8�}���Y���F�G1�*���#�1�<�
�>�}�JϮ�H¹��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��F���&����R��P �����&�{�x�_�w�}�(�������T9��D��*���6�o�%�:�2�.���UӖ��9��R	���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��9��h��\���=�;�_�u�w�}�W���Y����l��D��I���
�d�_�u�w�}�W������F�N��Uʥ�d�
�;�&�0�a�W���H����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�g�4��1�(���
����@��YN�����&�u�x�u�w�-�F݁�	����l��D�����2�
�'�6�m�-����
ۖ��9��h��Yʥ�d�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�*���#�1�|�!�2�}�W���Y���F��h_�����9�
�;�&�0�a�W���K����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�T��G1�����
�<�u�h�'�l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�g�>�����
������T��[���_�u�u�
�e�4�(���&����T��E��Oʥ�:�0�&�%�f�q���&����F��\�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`���&����_����ߊu�u�u�u�w�}�(�������TF���G�ߊu�u�u�u�;�8�}���Y���F�G1�*���&�2�i�u��o����B���F���U���u�u�u�0�3�-����
��ƹF��h_�����
�0�1�3��k�(��E���X��\�����2�u�!�0�$�c�Z���s���C9��R�����&�9�
�
��(�F��&����9l�N�U���`�4�
�9�w�.����	����@�CךU���
�`�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�`�;�(��M����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����%�6�;�!�;�l�G������\��h��D��
�g�|�|�#�8�W���Y���F���@���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�S��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�d�6���������l��^	�����u�u�'�6�$�u�(ށ�	����F��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ד�C9��SG�����u�u�u�u�w�}�WϮ�H����E
��^ �����h�%�d�4��1�L���Y�����RNךU���u�u�u�u����������@��S��*ۊ�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h�����4�&�2�u�%�>���T���F��1��*���
�&�<�;�'�2�W�������@N��B��*ۊ�'�2�u�
��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���#�1�|�!�2�}�W���Y���F��h_�����2�i�u�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�9�.���Y����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`�g�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L�֓�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����9�y�%�`�g�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�%�!�9���������h^�����1�_�u�u�w�}����s���F�N�����e�4�
�9��3����E�Ƽ�9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ƹ��Z��^	�����;�%�:�0�$�}�Z���YӖ��lV��Y1�����&�2�
�'�4�g��������lS��N��@���%�0�y�%�b�m������ƹF��R	�����u�u�u�3��<�(���
����T��N�����e�4�
�9�~�}����s���F�N�����e�<�
�<�w�`����I���F�N�����u�u�u�u�w�}����I����@��S��*ߊ�
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����V��G1�����
�<�u�&�>�3�������KǻN��*ߊ�e�4�
�9��3��������]9��X��U���6�&�}�
��m��������lS��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ӓ�9��h��\���=�;�_�u�w�}�W���Y����V��G1�����
�<�u�h�'�h�F߁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ӓ�9��h��*���&�2�i�u���G���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`�f�����Ӈ��Z��G�����u�x�u�u�'�h�F߁�����l��^	�����u�u�'�6�$�u�(ځ�I�Ƽ�9��h�����
�
�e�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�*���#�1�|�!�2�}�W���Y���F��h[��E���
�<�u�h�'�h�F��Y���F��[�����u�u�u�u�w��(�������TF���*���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�9��h��*���&�2�4�&�0�}����
���l�N��@��
�%�#�1�>�����
����l��TN����0�&�%�`�f������Ƽ�9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ƹ��l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�9��h��*���&�2�i�u���F���&����9F�N��U���0�_�u�u�w�}�W���&ƹ��l��A�����<�u�h�%�b�l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�f�4�(���Y����T��E�����x�_�u�u���F���&����R��P �����o�%�:�0�$�-�B��UӖ��lW��G��Yʥ�`�d�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h_�����9�|�u�=�9�W�W���Y���F��1�*���&�2�i�u���F�ԜY���F��D��U���u�u�u�u�'�h�Fށ�����Z�G1��Dۊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ƹ��l��A�����<�u�&�<�9�-����
���9F���*���4�
�9�
�9�.����
����C��T�����&�}�
�
�e�<�(���UӖ��lW��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�L����R��[
��U���;�_�u�u�w�}�W���&ƹ��l��A�����<�u�h�%�b�l�(�������F�N�����u�u�u�u�w�}�WϮ�L����R��[
�����2�i�u�
��o��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�`�d��3��������]F��X�����x�u�u�%�b�l�(���
����@��Y1�����u�'�6�&���(��Y����T��E��U���
�g�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��\�����1�|�!�0�w�}�W���Y�����h_�����<�u�h�%�b�l�L���Y�����RNךU���u�u�u�u���E���&����[��h[��G���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�L����R��[
�����2�4�&�2�w�/����W���F�G1��Dي�%�#�1�<��4�(�������A	��N�����&�%�`�d��-����Y����U��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&�Փ�C9��SG�����u�u�u�u�w�}�WϮ�L����R��[
�����2�i�u�
��n������ƹF�N�����_�u�u�u�w�}�W���&�Փ�C9��S1��*���u�h�%�`�f���������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�f�>�����
������T��[���_�u�u�
��n��������@��h����%�:�0�&�'�h�F��	�ӓ� 9��R	����d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lS��1��*���|�u�=�;�]�}�W���Y���C9��]�����2�i�u�
��n�}���Y���V
��d��U���u�u�u�%�b�l�(���
���F��1�*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&�ғ�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h[��A���
�9�
�;�$�:��������\������}�
�
�a�6����	�ӓ�9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����Hǹ��l��G�����_�u�u�u�w�}�W���&�ғ�C9��S1��*���u�h�%�`�f��������F�N�����u�u�u�u�w�}����Hǹ��l��h�����i�u�
�
�c�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�`�d�
�9�.�Ͽ�
����C��R��U���u�u�%�`�f���������Z��G��U���'�6�&�}���C���&ƹ��l��PB��*ߊ�a�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��h�����|�!�0�u�w�}�W���Y����lS��1��*���u�h�%�`�f�f�W���Y����_��=N��U���u�u�u�
��i���������h_�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����Hƹ��l��h�����4�&�2�u�%�>���T���F��1�*���#�1�<�
�>���������PF��G�����%�`�d�
�'�+����&ƹ��l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ځ�L����E
��N�����u�u�u�u�w�}����Hƹ��l��h�����i�u�
�
�b�<�(���B���F����ߊu�u�u�u�w�}�(ځ�L����E
��^ �����h�%�`�d��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�`�<��4�W�������A	��D�X�ߊu�u�
�
�b�4�(���&����T��E��Oʥ�:�0�&�%�b�l�[Ϯ�L����C��N��@��
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lW��V�����u�=�;�_�w�}�W���Y�Ƽ�9��h�����i�u�
�
�b�W�W���Y�Ʃ�@�N��U���u�u�%�`�f��������C9��[�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ځ�&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�;�&�2�6�.���������T��]���
�
�%�#�3�}�(ځ�&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�b�l�������G��d��U���u�u�u�%�b�l��������l��R�����d�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
��-��������TF���*ۊ�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h_�����2�4�&�2�w�/����W���F�G1��D���
�<�
�&�>�3����Y�Ƽ�\��DF��@��u�
�
�
�%�:�W���&¹��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��-����PӒ��]FǻN��U���u�u�
�
��3����E�Ƽ�9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��^ �����h�%�`�d�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h[��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
�'�+����&����R��P �����o�%�:�0�$�-�B�������WJ��h[��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��V�����;�&�2�i�w��(݁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ӓ�l��A�����<�u�h�%�b�o��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�`�g�>�����
������T��[���_�u�u�
����������Z��G��U���'�6�&�}���[Ϯ�L�ԓ�A����*؊�%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ӓ�l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�l��D��I���
�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�;�$�:�K���&ƹ��C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`�d�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L�Փ�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����9�y�%�`�d�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�%�!�9���������h]�����1�_�u�u�w�}����s���F�N�����f�4�
�9��3����E�Ƽ�9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ƹ��Z��^	�����;�%�:�0�$�}�Z���YӖ��lU��Y1�����&�2�
�'�4�g��������lS��N��@���%�0�y�%�b�n������ƹF��R	�����u�u�u�3��<�(���
����T��N�����f�4�
�9�~�}����s���F�N�����f�<�
�<�w�`����J���F�N�����u�u�u�u�w�}����J����@��S��*ߊ�
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��h��*���&�2�4�&�0�}����
���l�N��@���4�
�9�
�9�.����
����C��T�����&�}�
�
��-����Y����9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����M����E
��N�����u�u�u�u�w�}����M����E
��^ �����h�%�`�a�6����Y���F��[�����u�u�u�u�w��(ہ�	����l��D��I���
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�
�;�&�2�6�.��������@H�d��Uʥ�`�a�<�
�>���������PF��G�����%�`�a�u���(����Ƽ�9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(ہ�	����O��_�����u�u�u�u�w��(ہ�����Z�G1��A�ߊu�u�u�u�;�8�}���Y���F�G1��A���
�<�u�h�'�h�C�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(�������]9��P1�����
�'�6�o�'�2����	�ӓ�l��A��U���
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��@���
�9�|�u�?�3�}���Y���F�G1��@���
�9�
�;�$�:�K���&ƹ��R��[
�U���u�u�0�&�w�}�W���Y�����h[�����1�<�
�<�w�`����L����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h�B���&����R��P �����&�{�x�_�w�}�(ځ�&����Z��D�����:�u�u�'�4�.�_���&����lS��h�����
�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h[�����1�|�!�0�w�}�W���Y�����h[�����2�i�u�
��f�W���Y����_��=N��U���u�u�u�
���������C9��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�B�������W9��h��U���<�;�%�:�2�.�W��Y����lS��h�����<�
�<�
�$�4��������C��R�����c�4�
�9�{�-�B�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
����������[��=N��U���u�u�u�
����������@��S��*ߊ�
�%�#�1�]�}�W���Y����l�N��U���u�%�`�c�6���������Z�G1��C���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��1��*���u�&�<�;�'�2����Y��ƹF��h[��*���&�2�4�&�0�����CӖ��P����*���%�`�c�%�2�q����O����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�`�c�6�����Y����l�N��U���u�%�`�c�>�����DӖ��lP��N��U���0�&�u�u�w�}�W���YӖ��lP��Y1����u�
�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�����9�
�;�&�0�<����Y����V��C�U���%�`�b�4��1�(���
����@��Y1�����u�'�6�&���(؁�	����F��1�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lQ��G1�����!�0�u�u�w�}�W���YӖ��lQ��G1�����
�<�u�h�'�h�@���&����9F�N��U���0�_�u�u�w�}�W���&ƹ��R��[
�����2�i�u�
����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
�9�.�Ͽ�
����C��R��U���u�u�%�`�`�4�(���&����T��E��Oʥ�:�0�&�%�b�j�W���&Ĺ��V�G1��B���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ƹ��R��[
��U���;�_�u�u�w�}�W���&ƹ��Z��^	��Hʥ�`�b�_�u�w�}�W������F�N��Uʥ�`�b�<�
�>�}�JϮ�L�ѓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&˹��l��h�����4�&�2�
�%�>�MϮ�������hV�����1�u�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�`�m�4�
�;�t�W������F�N��Uʥ�`�m�4�
�;��������C9��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�
�%�#�1�>�����DӖ��l^��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�L�ޓ�]9��PN�����u�'�6�&�y�p�}���Y����9��h��*���<�;�%�:�w�}����
�μ�9����*Ҋ�'�2�u�
���������F��P��U���u�u�<�u��-��������Z��S��*ߊ�
�%�#�1�~�)����Y���F�N��*ߊ�
�;�&�2�k�}�(ځ�B���F����ߊu�u�u�u�w�}�(ځ�&����Z�
N��@���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�l��A�����<�u�&�<�9�-����
���9F���*ӊ�%�#�1�<��4�(�������A	��N�����&�%�`�l�6����	�ӓ�l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ځ�&����_����ߊu�u�u�u�w�}�(ځ�&����_��Y1����u�
�
�
�'�+��ԜY���F��D��U���u�u�u�u�'�h�N���&����Z��^	��Hʥ�`�l�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��@���<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�;�&�0�<����&����\��E�����
�
�y�%�b�d����UӖ��l_��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�h�N���&����F��R ��U���u�u�u�u�'�h�N���&����[��h[��N���u�u�u�0�$�}�W���Y���F��h[��*���&�2�i�u���(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����e�4�
�9��3��������]F��X�����x�u�u�%�`�m��������l��h�����%�:�u�u�%�>����&Ĺ��R��[
����e�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*���#�1�|�!�2�}�W���Y���F��hY��*���#�1�<�
�>�}�JϮ�N�֓�C9��SUךU���u�u�9�0�]�}�W���Y���C9��1��*���
�;�&�2�k�}�(؁�&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(���
����@��YN�����&�u�x�u�w�-�@�������T9��D��*���6�o�%�:�2�.����I�Ƽ�9��G��Yʥ�b�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��1��*���|�u�=�;�]�}�W���Y���C9��1��*���u�h�%�b�g�W�W���Y�Ʃ�@�N��U���u�u�%�b�g�4�(���Y����lQ��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������W9��h��U���<�;�%�:�2�.�W��Y����lQ��1��*���
�;�&�2�6�.���������T��]���
�e�4�
�;�q����Hù��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�j�F߁�	����O��_�����u�u�u�u�w��(�������W9��h��U��%�b�d�
�'�+��ԜY���F��D��U���u�u�u�u�'�j�F߁�	����l��D��I���
�
�e�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����d�
�;�&�0�<����Y����V��C�U���%�b�d�
�9�.����
����C��T�����&�}�
�
�g�}�(؁�I����TJ��hY��E���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��l��A��\ʡ�0�u�u�u�w�}�W���	�ѓ�9��h��U��%�b�d�n�w�}�W�������9F�N��U���u�
�
�e�>�����DӖ��lW��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�Fށ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��h�����<�
�<�
�$�4��������C��R�����d�
�%�#�3�}�(؁�H����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���F���&����F��R ��U���u�u�u�u�'�j�Fށ�	����l��D��I���
�
�d�4��1�L���Y�����RNךU���u�u�u�u���F���&����Z��^	��Hʥ�b�d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�d�<�
�<�w�.����	����@�CךU���
�
�d�<��4�(�������A	��N�����&�%�b�d�{�-�@��&����F�� 1�*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�N����R��[
��U���;�_�u�u�w�}�W���&Ĺ��l��D��I���
�
�d�_�w�}�W������F�N��U���%�b�d�
�9�.���Y����W��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���E���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��lW��V�����;�&�2�4�$�:�(�������A	��D��*݊�g�4�
�9�{�-�@��&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`�l�(��������YNךU���u�u�u�u���E���&����Z��^	��Hʥ�b�d�
�%�!�9�}���Y���V
��d��U���u�u�u�%�`�l�(�������]9��PN�U���
�g�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B��
�;�&�2�6�.��������@H�d��Uʥ�b�d�
�;�$�:��������\������}�
�
�g�w��(���	������h_�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&�ԓ�C9��SG�����u�u�u�u�w�}�WϮ�N����Z��^	��Hʥ�b�d�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�g�<��4�W��	�ѓ�9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`�l�(�������]9��PN�����u�'�6�&�y�p�}���Y����U��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B��
�%�#�1�w��(�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��n�������G��d��U���u�u�u�%�`�l�(�������]9��PN�U���
�f�4�
�;�f�W���Y����_��=N��U���u�u�u�
��n��������l��R�����d�
�%�#�3�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�f�<�
�>���������PF��G�����%�b�d�y�'�j�F܁����C9��]�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����H����l��G�����_�u�u�u�w�}�W���&�Փ�]9��PN�U���
�f�_�u�w�}�W������F�N��Uʥ�b�d�
�;�$�:�K���&Ĺ��l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��i��������l�������%�:�0�&�w�p�W���	�ѓ�9��h��*���&�2�4�&�0�����CӖ��P����*���4�
�9�y�'�j�Fہ�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�b�f���������[��=N��U���u�u�u�
��i��������l��R�����d�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�b�f���������@��S��*݊�a�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��Dފ�;�&�2�4�$�:�W�������K��N�����d�
�;�&�0�<����&����\��E�����
�
�a�u���C�������lQ��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(؁�M����E
��N�����u�u�u�u�w�}����Hǹ��l��R�����d�n�u�u�w�}����Y���F�N��U���
�a�<�
�>�}�JϮ�N����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b�f���������@��V�����'�6�&�{�z�W�W���&Ĺ��l��A�����<�
�&�<�9�-����Y����V��G1��Dߊ�%�#�1�u���B���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�b�<�(���P�Ƹ�V�N��U���u�u�%�b�f���������@��S��*݊�`�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
�b�<�(���&����Z�
N��B��
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��@���
�<�u�&�>�3�������KǻN��*݊�`�<�
�<��.����	����	F��X��¥�b�d�y�%�`�l�(����Ƽ�9��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@��&����_����ߊu�u�u�u�w�}�(؁�L����@��S��*݊�`�_�u�u�w�}����s���F�N�����d�
�;�&�0�a�W���&�ӓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&¹��l��h�����4�&�2�
�%�>�MϮ�������h_�����1�u�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b�d�4�
�;�t�W������F�N��Uʥ�b�d�4�
�;��������C9��1��*���n�u�u�u�w�8����Y���F�N��*݊�
�%�#�1�>�����DӖ��lW��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�N�ד�]9��PN�����u�'�6�&�y�p�}���Y����9��h��*���<�;�%�:�w�}����
�μ�9����*ۊ�'�2�u�
���������F��P��U���u�u�<�u��-��������Z��S��*݊�
�%�#�1�~�)����Y���F�N��*݊�
�;�&�2�k�}�(؁�B���F����ߊu�u�u�u�w�}�(؁�&����Z�
N��B���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�l��A�����<�u�&�<�9�-����
���9F���*؊�%�#�1�<��4�(�������A	��N�����&�%�b�g�6����	�ѓ�l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(؁�&����_����ߊu�u�u�u�w�}�(؁�&����_��Y1����u�
�
�
�'�+��ԜY���F��D��U���u�u�u�u�'�j�E���&����Z��^	��Hʥ�b�g�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�;�&�0�<����&����\��E�����
�
�y�%�`�o����UӖ��lT��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�j�E���&����F��R ��U���u�u�u�u�'�j�E���&����[��hY��N���u�u�u�0�$�}�W���Y���F��hY��*���&�2�i�u���(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����f�4�
�9��3��������]F��X�����x�u�u�%�`�n��������l��h�����%�:�u�u�%�>����&Ĺ��R��[
����f�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*���#�1�|�!�2�}�W���Y���F��hY��*���#�1�<�
�>�}�JϮ�N�Փ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��1��*���
�;�&�2�k�}�(؁�&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(���
����@��YN�����&�u�x�u�w�-�@�������T9��D��*���6�o�%�:�2�.����J�Ƽ�9��G��Yʥ�b�f�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��1��*���|�u�=�;�]�}�W���Y���C9��1��*���u�h�%�b�d�W�W���Y�Ʃ�@�N��U���u�u�%�b�d�4�(���Y����lQ��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(ہ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��V�����;�&�2�4�$�:�(�������A	��D��*݊�
�%�#�1�w��(ہ�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�b�c�<�(���P�Ƹ�V�N��U���u�u�%�b�c�<�(���&����Z�
N��B���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
�'�+����&����[��hY��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lQ��h�����4�&�2�u�%�>���T���F�� 1�����<�
�&�<�9�-����Y����V��G1��A���
�
�
�'�0�}�(؁�&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�'�+��������9F�N��U���u�
�
�
�9�.���Y����]ǻN��U���9�0�_�u�w�}�W���Y����9��h��U��%�b�a�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h[�����1�<�
�<�w�.����	����@�CךU���
�
�
�%�!�9��������@��h����%�:�0�&�'�j�B���&������h[�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����9��h��\���=�;�_�u�w�}�W���Y����9��h��*���&�2�i�u���(�������F�N�����u�u�u�u�w�}�WϮ�N�ӓ�C9��S1��*���u�h�%�b�b�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b�`�<��4�W�������A	��D�X�ߊu�u�
�
��3��������]9��X��U���6�&�}�
��q����L����TJ��hY��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�N�ӓ�C9��SG�����u�u�u�u�w�}�WϮ�N�ӓ�]9��PN�U���
�n�u�u�w�}����Y���F�N��U���
�
�;�&�0�a�W���&ƹ��V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�b�c�6�����������^	�����0�&�u�x�w�}����O����E
��^ �����&�<�;�%�8�}�W�������C9��1��*���y�%�b�c�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�%�#�3�t����Y���F�N��U���
�
�%�#�3�4�(���Y����lQ��h�����_�u�u�u�w�1��ԜY���F�N��B���4�
�9�
�9�.���Y����9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&Ź��l�������%�:�0�&�w�p�W���	�ѓ�l��D�����2�
�'�6�m�-����
ۖ��lP�G1��C���0�y�%�b�a�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��B���4�
�9�|�w�5��ԜY���F�N��B���<�
�<�u�j�-�@��s���F�R��U���u�u�u�u�w�-�@�������TF���*܊�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&Ĺ��R��[
�����2�4�&�2�w�/����W���F�G1��B���
�9�
�;�$�:��������\������}�
�
�
�'�+����&Ĺ��R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@�������WO�C��U���u�u�u�u�w�-�@�������W9��h��U��%�b�b�4��1�L���Y�����RNךU���u�u�u�u���(�������]9��PN�U���
�
�%�#�3�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*݊�;�&�2�4�$�:�W�������K��N�����b�<�
�<��.����	����	F��X��¥�b�b�u�
������Y����9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(��������YNךU���u�u�u�u���(���
���F�� 1����u�u�u�9�2�W�W���Y���F�� 1�����<�u�h�%�`�j����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�%�#�1�>�����
������T��[���_�u�u�
����������@��V�����'�6�o�%�8�8�Ǯ�N�ޓ�C9��SB��*݊�
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F�� 1�����9�|�u�=�9�W�W���Y���F�� 1�����9�
�;�&�0�a�W���&˹��l��d��U���u�0�&�u�w�}�W���Y����lQ��h�����<�
�<�u�j�-�@�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`�e�����ƭ�@�������{�x�_�u�w��(ׁ�����l��^	�����u�u�'�6�$�u�(؁�UӖ��l^��E��U���
�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lQ��h�����|�!�0�u�w�}�W���Y����lQ��h�����i�u�
�
�l�}�W���YӃ��VFǻN��U���u�u�
�
��3����E�Ƽ�9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�N���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l_��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B���4�
�9�y�'�j�N���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��-����PӒ��]FǻN��U���u�u�
�
��-��������TF���*ӊ�%�#�1�_�w�}�W������F�N��U���%�b�l�4��1�(���
���F�� 1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��^ �����&�<�;�%�8�8����T�����hW�����2�4�&�2��/���	����@��hY��Yʥ�b�l�%�0�{�-�@�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b�l�4��1�^������F�N��U���%�b�l�<��4�W��	�ѓ�l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�l��D��I���
�
�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����[�I�����}�8�
�
�"�l�Eׁ�K����C9��Y����
�|�0�&�w�l�L�ԜY�����h�����4�&�2�u�%�>���T���F��1��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������F��^�����3�
�d�a�'�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Y������T�����d�e�h�0�>�>��������R��G��\ʡ�0�u�u�u�w�}�W���	�ޓ�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�e���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����R��[
�����2�4�&�2�w�/����W���F�G1�����9�
�;�&�0�<����&����\��E�����
�
�%�#�3�}�(ց�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l�6�����Y����l�N��U���u�%�l�4��1�(���
���F��1��*���n�u�u�u�w�8����Y���F�N��*ӊ�%�#�1�<��4�W��	�ߓ�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�N���&����R��P �����&�{�x�_�w�}�(ց�����l��^	�����u�u�'�6�$�u�(��	�ߓ�A����*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�@����E
��N�����u�u�u�u�w�}��������TF���N���u�u�u�0�$�}�W���Y���F��hW�����2�i�u�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��D��*ߊ�
� �d�`��l�W��Q���N�F��]´�'�9�
�:��2���&�ӓ�9��h\�U���'�
�!��%�����N����R��B1�M���u�'�
�!��/�;���&�ѓ�9��h��G��u�u�'�
�#���������lW��\�� ��e�u�u�'��)�1���5����Q��1�*���g�c�u�u�%���������C9��h_��Dڊ� �g�g�u�w�/�(���?����\	��Y��@���3�
�c�|�q�<����&����	��h\��Dߊ�
� �g�a�w�}��������l*��G1�*���b�3�
�c�~�{��������A9��X��B��
�
� �g�a�}�W���&����\��X��G݊�`�`�3�
�b�t�QϿ�����u	��{��*���d�
�
� �e�e�W�������l ��h"����
�`�f�3��i�^�������G9��E1�����b�d�
�
�"�o�G���Y����_��X�����g�
�`�d�1��D���_Ӈ��l
��q��9���
�b�d�
�"�o�E��Y����l4��B��C���3�
�`�d�'�j�K���Q���N�F��]���
�!��'��2�(���Hƹ��l ��[�Sʴ�'�9�
�:��2���&�ӓ�9��h]�\��4�'�9�
�8�����Kʹ��lW��Q��A���s�4�'�9��2�(���	����S��1��*��|�s�4�'�;���������
9��h_�����a�|�s�4�%�1�(���&����lT��[��E���
�f�|�s�6�/��������\��1�*ӊ� �f�g�u�w�/�(���?����\	��W��@���3�
�g�|�q�<����&����	��h\��Dߊ�
� �f�a�w�}��������l*��G1�*���c�3�
�g�~�{��������A9��X��L��
�
� �f�a�}�W���&����\��X��Gӊ�`�a�3�
�f�t�QϿ�����u	��{��*���d�
�
� �d�e�W�������l ��h"����
�`�g�3��m�^�������G9��E1�����l�d�
�
�"�n�G���Y����_��X�����g�
�`�3��d�^�ԜY�Ƹ�C9��h_�C���u�h�<�
�>���������A��W�A���d�1�"�!�w�t�}���Y����@9��h_�M���u�h�}�
�2�(����
����S��h�U���%��&�9���(���H����CW��d��Uʠ�
����"��N���&����CU�
NךU���u�u�%�6�9�)���&�ƻ�V�U��*���,� �
�b�1��Cہ�K���F�G�����_�u�u�u�w��F���&����9������