-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��l��e��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e��"��g�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӇ��P�'��&������_�w�}�(߁�����9��h��U���������}���Y����a��~1�Oʜ�u��
����2���+������Y��E��u�u�%�e��*�>�������WF��~ ��!�����n�u�w�-�G�������\��yN��1��������}�F�������V�=N��U���
�4��
��-����Cӯ��`2��{!��6�ߊu�u�
�
�6��(���Y����g"��x)��*�����}�`�3�*����P���F��1�����f�4�
�9�w�}�9ύ�=����z%��N������"��a�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�֓�R��hZ�����1�o��u���8���B�����h<��4���u�u�����0���/����aF�N�����u�|�_�u�w��(���8����R��[
��U��������W�W���&ù��D'��N�<����
�����#���Q����\��XN�N���u�%�e�� ��A���&����	F��=��*����n�u�u�'�m�%���0���/��d:��9�������w�l�W������]ǻN��*ڊ�4��
�
�'�+���0�Ɵ�w9��p'�����u�
�
�4���W���7ӵ��l*��~-��0����}�`�1� �)�W���s���C9��e��<���4�
�9�u�w��$���5����l�N��E���"��l�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I����r/��h�����o��u����>��Y����lV��V��*��o��u����>���<����N��
�����e�n�u�u�'�m�%���0����R��[
��U��������W�W���&ù��D'��_��U���������4���Y����W	��C��\�ߊu�u�
�
�6��(�������WF��~ ��!�����n�u�w�-�G�������F��~ ��!�����
����_������\F��d��Uʥ�e��"��f���������}F��s1��2���_�u�u�
��<�6���J����}F��s1��2������u�f�}�������9F���*����
�f�4��1�W���7ӵ��l*��~-�U���%�e��"��l�W���7ӵ��l*��~-��0����}�`�1� �)�W���s���C9��e��<��
�%�#�1�m��W���&����p]ǻN��*ڊ�4��
�`�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�֓�R��h_�����9�u�u����;���:���F��1������
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�M����_��~1�����9�u�u� �w�	�(���0��ƹF��hZ�����1��d�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ǹ��R
��v'��*���#�1�o����3���>����F�G1��&���0��
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ғ�P��S/��G���
�9�u�u��}�#���6����9F���*���9�1��f�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����`��R
��*ي�%�#�1�o��	�$���5����l�N��A���4�0��
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l5��[��<���4�
�9�u�w��W���&����p]ǻN��*ފ�6�9�1��b�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�9��V��4���
�%�#�1�m��#ύ�=����z%��N������4�0���}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lR��T�����c�4�
�9�w�}�"���-����t/��=N��U���
�6�9�1��j�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���C9��d�����
�
�%�#�3�g�8���*����|!��d��Uʥ�a��4�0���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h=������m�4�
�;�}�W���Y����)��tUךU���
�
�6�9�3��N��6����g"��x)��*�����}�d�3�*����P���F��1������
�
�%�!�9�Mϑ�-ӵ��l*��~-�U���%�a��4�2��(��Cө��5��h"��<������}�f�9� ���Y����F�G1��&���0��
�e�6�����Y����`2��{!��6�ߊu�u�
�
�4�1����H����|3��d:��9�������w�n�W������]ǻN��*ފ�6�9�1��f���������f2��c*��:���n�u�u�%�c�����8����\��b:��!�����
����_������\F��d��Uʥ�a��4�0���E���&����	F��cN��1�����_�u�w��(�������lW��N��!ʆ�������8���J�ƨ�D��^����u�
�
�6�;�9�>��&����_�!��U���
���n�w�}����*����W'��Z��U���u��
����2���+������Y��E��u�u�%�a��<����&�ғ�C9��SN�:��������W�W���&ǹ��R
��v'��@��������4���:����U��S�����|�_�u�u����������9��h��U��� �u��
���L���YӖ��l$��T��;ʆ�������8���H�ƨ�D��^����u�
�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��1��*���u�u�����0���s���C9��u1�Oʜ�u��
����2���+������Y��E��u�u�%�b��o��������z(��c*��:���n�u�u�%�`��D��0�Ɵ�w9��p'��#����u�d�u�8�3���B�����h,��*���#�1�o��w�	�(���0��ƹF��hY��*���u������4���:����W��S�����|�_�u�u���(ہ�	����\��yN��1�����_�u�w��(���Y�ƅ�5��h"��<������}�b�9� ���Y����F�G1��7���4�
�9�u�w��$���5����l�N��B���c�o��u���8���&����|4�[�����:�e�n�u�w�-�@���O����E
��N��U���
���n�w�}����;���/��d:��9�������w�l�W������]ǻN��*݊�
�
�%�#�3�g�>���-����t/��=N��U���
�
�u�u���3���>����v%��eN��@ʱ�"�!�u�|�]�}�W���&����R��[
��U��������W�W���&Ĺ��
F��~ ��!�����
����_������\F��d��Uʥ�b��l�4��1�W���7ӵ��l*��~-�U���%�b��d�w�}�9ύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����q9��h�����o��u����>��Y����lQ��h_�Oʜ�u��
����2���+������Y��E��u�u�%�b��l�(������/��d:��9����_�u�u���(��Cӯ��`2��{!��6�����u�d�w�2����I��ƹF��hY��*���4�
�9�u�w��$���5����l�N��B���d�u�u����;���:����g)��_����!�u�|�_�w�}�(؁�&�Փ�C9��SN�<����
���l�}�WϮ�N����F��~ ��!�����
����_������\F��d��Uʥ�b��d�
�'�+���0�Ɵ�w9��p'�����u�
�
�
�b�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӖ��l$��1��*���u�u�����0���s���C9��z1�Oʜ�u��
����2���+������Y��E��u�u�%�l��m��������z(��c*��:���n�u�u�%�n��F��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h#��*���#�1�o��w�	�(���0��ƹF��hW��*���u������4���:����U��S�����|�_�u�u���(݁�	����\��yN��1�����_�u�w��(���Y�ƅ�5��h"��<������}�f�9� ���Y����F�G1��8���4�
�9�u�w��$���5����l�N��L���a�o��u���8���&����|4�_�����:�e�n�u�w�-�N���M����E
��N��U���
���n�w�}����4���/��d:��9�������w�n�W������]ǻN��*ӊ�
�
�%�#�3�g�>���-����t/��=N��U���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����R��[
��U��������W�W���&ʹ��F��~ ��!�����
����_������\F��d��Uʥ�l��b�4��1�W���7ӵ��l*��~-�U���%�l��m�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ߓ�l^��G1�����u��
���L���YӖ��l+��T��;ʆ�������8���J�ƨ�D��^����u�
�
�
��-����Cӯ��`2��{!��6�ߊu�u�
�
��m�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����l_��h_�����9�u�u����;���:���F��1��D���u������4���:����U��S�����|�_�u�u���(�������WF��~ ��!�����n�u�w�-�N���H����z(��c*��:���
�����l��������l�N��L���d�
�%�#�3�g�>���-����t/��=N��U���
�
�f�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�@���� 9��h��U���������}���Y����~9��T��;ʆ�������8���J�ƨ�D��^����u�
�
�
�c�<�(���Y�ƅ�5��h"��<��u�u�%�l��l�W���7ӵ��l*��~-��0����}�d�1� �)�W���s���C9��z1�*���#�1�o��w�	�(���0���9��dװ���<�0�!�'�w�8����Ӌ��_��^��Eʼ�u�u�u�4�#�4����:����t#��e/��:�����o����L���YӇ��A��C��:���������9����Ʈ�[��N�����0�!�'�u�$�}�W���L����wW��h^�����%�g�d�
�{��$���)����j6��T��=��������	�FÖ�*����f2��~6��H����
�� ���#Ҧ�N����P
��Z��Y���
�� �
���J��I����J��d1��%�����h�!�2�.�?���*����)��
_�L��e�y��
���6��@߮��l5��h:��H���0������:��1����j(��d>��Y���
��
��f�m�[���&����3��W���u�u�6�;�#�3�W�������l
��^��U����
���w�`�P���s���P	��C��U���6�;�!�9�0�>�G��*����|!��T��R��_�u�u�:�$�<�Ͽ�&����GW��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��B�����D��ʴ�
��&�g�1�0�F��*����|!��h8��!���}�f�1�"�#�}�^��Y����V��^�E��n�u�u�6�9�)����	����@��Q��G��������4���Y����W	��C��\��u�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�D��w�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�F��I��ƹF��X �����4�
��&�a�;���Cӵ��l*��~-��0����}�f�1� �)�W���C���V��^�E��e�n�u�u�4�3����Y����g9�� 1����o������!���6��� F��@ ��U���o�u�e�e�g�m�G��I����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�w�_�u�w�2����Ӈ��`2��CW�����u�u��
���(���-���U��X����u�h�w�e�g�l�G��I���9F������!�4�
��$�l�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�e�w�_�w�}��������C9��h��D���8�d�u�u���8���&����|4�]�����:�e�u�h�u�m�F��I����V�=N��U���&�4�!�4��	���&����W�=��*����
����u�DϺ�����O�
N��E��e�e�e�e�g�f�W�������R��V��!���d�
�&�
�e�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�N���u�6�;�!�9�}����&����l ��h_�Oʆ�������8���H�ƨ�D��^��O���d�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�F��*����|!��h8��!���}�u�:�;�8�m�W��[����F�T�����u�%�6�;�#�1�Fف�Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����d�e�o����0���/����aF�
�����e�u�h�w�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������qF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�D��u�u�6�;�#�3�W�������l
��h^��U���
���
��	�%���Y����G	�N�U��e�e�n�u�w�>�����ƭ�l��D�����e�o�����4���:����P��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�d�n�w�}��������R��X ��*���a�g�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����c�
�u�u���8���&����|4�]�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�a�a�o���;���:����g)��X����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�c�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�d�f�f�W�������R��V�����
�#�a�c�m��3���>����v%��eN��Fʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�c�
�w�}�#���6����e#��x<��C���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�f�l�L���YӅ��@��CN��*���&�
�#�a�o�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�c��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�F��Y����\��V �����:�&�
�#�c��Mύ�=����z%��r-��'���f�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�l�F���s���P	��C��U���6�;�!�9�a��W���-����t/��a+��:���c�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�i�4��*����|!��h8��!���}�f�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�k�(���Y����)��t1��6���u�c�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��H��ƹF��X �����4�
�:�&��+�C���Cӵ��l*��~-��0����}�f�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�Aہ�Y�Ɵ�w9��p'��#����u�c�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��H���9F������!�4�
�:�$�����=����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���&���5��h"��<������}�w�2����I����D��^�N���u�6�;�!�9�}��������ER��T��!�����
����_�������V�S��E��w�_�u�u�8�.��������]��[��A��������4���Y����\��XN�U��w�d�e�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�f��}���Y����G�������!�9�a�m�m��3���>����v%��eN��U���;�:�e�u�j��G��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���f�1�"�!�w�t�M���H����l�N�����;�u�%�6�9�)����:����g"��x)��*�����}�u�8�3���Y���W��UךU���:�&�4�!�6�����&����F��d:��9�������w�n��������\�^�E��u�u�6�;�#�3�W�������l
��h_��U���
���
��	�%���Y����G	�N�U��e�w�_�u�w�2����Ӈ��P	��C1��A��o������!���6�����Y��E���h�w�e�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�U�ԜY�Ư�]��Y�����;�!�9�a�`�g�$���5����l0��c!��]���:�;�:�e�w�`�U��H��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�f�1�"�#�}�^��Y����D��N�����!�;�u�%�4�3����M���5��h"��<������}�w�2����I����D��_�����u�:�&�4�#�<�(���
����9��N��1��������}�DϺ�����O�
N��D��n�u�u�6�9�)����	����@��A[��U����
�����#���Q�ƨ�D��^��O���e�e�e�n�]�}�W�������C9��h��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��B�����E�����&�
�;�:�>�:�Mϭ�����9F������!�u�&�
�9�2�����ƭ�l%��Q��Oʦ�2�4�u�&�u�2���Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&���� V�,��9���n�u�u�&�0�<�W���&����z9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(߁�����9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"��e�6���������\��c*��:���n�u�u�&�0�<�W���&����z9��V�����'�2�o����0���C���]ǻN�����9�%�e�� ��F���&����	F��s1��2������u�f�}�������9F������%�e��"��l����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l4��v'��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�e�� ��F���&����C��T��!�����u�h�p�z�}���Y����R
��h^�����
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h<��4���
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u������&����l��h�����o������}���Y����R
��h^�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����z9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(߁����� 9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"��f�6���������\��c*��:���n�u�u�&�0�<�W���&����z9��V�����'�2�o����0���C���]ǻN�����9�%�e�� ��C���&����	F��s1��2������u�f�}�������9F������%�e��"��i����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l4��v'��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�e�� ��C���&����C��T��!�����u�h�p�z�}���Y����R
��h^�����
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h<��4���
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u������&ƹ��l��h�����o������}���Y����R
��h^�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����z9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(߁�����9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"��c�6���������\��c*��:���n�u�u�&�0�<�W���&����z9��V�����'�2�o����0���C���]ǻN�����9�%�e�� ��@���&����	F��s1��2������u�f�}�������9F������%�e��"��j����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l4��v'��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�e�� ��@���&����C��T��!�����u�h�p�z�}���Y����R
��h^�����
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h<��4���
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u������&˹��l��h�����o������}���Y����R
��h^�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����z9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(߁�����
9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"��l�6���������\��c*��:���n�u�u�&�0�<�W���&����z9��V�����'�2�o����0���C���]ǻN�����9�%�e�� ��F߁�����\��c*��:���
�����h��������l�N�����u�
�
�4���G�������`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�w�]�}�W�������lV��V��*���4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
��<�6���I����E
��G��U����
���w�`�P���s���@��V��*ڊ�4��
�d�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��E���"��d�
�%�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�M���I����V��^�E��n�u�u�&�0�<�W���&����z9��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�e��"��f���������TF��d:��9����o�u�e�l�}�Wϭ�����C9��e��<��
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lV��V��*���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�g�� ���H����l��h�����o������}���Y����R
��h^�����
�g�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�I����r/��1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&����z9��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�4���n��������l��T��!�����n�u�w�.����Y����a��~1�*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u������&�ғ�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�g�� ���Hǹ��V�=��*����
����u�BϺ�����O�
N��E��e�e�e�e�g�m�L���Yӕ��]��G1��'����d�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G�������9��h��*���2�o�����4��Y���9F������%�e��"��l�(���
���5��h"��<������}�b�9� ���Y����F�D�����
�
�4���h����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l4��v'��@���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�6��(�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lQ��h^�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�N����l��A�����u�u��
���W��^����F�D�����
�
�
�
�9�.���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T����*���
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u���(ށ�	����l��D��Oʆ�����]�}�W�������lQ��h_�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
���(���
���5��h"��<������}�b�9� ���Y����F�D�����
�
�
�
�%�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�M���I����V��^�E��n�u�u�&�0�<�W���&����R��[
�����2�o�����4�ԜY�ƿ�T����*���
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(؁�&����l��T��!�����
����_������\F��d��Uʦ�2�4�u�
���(�������g"��x)��*�����}�`�3�*����P���V��^�E��e�e�e�n�w�}�����Ƽ�9��1��*���
�;�&�2�m��3���>����F�D�����
�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����q9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(؁�&ǹ��V�=��*����
����u�BϺ�����O�
N��E��e�e�e�e�g�m�L���Yӕ��]��G1��7���4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
���(�������A��N��1�����o�u�g�f�W���
����_F�� 1��@���
�<�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����q9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�b��`�4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�&ƹ��l��h���������g�W��B�����Y������c�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F�� 1��C���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b��k��������l��T��!�����n�u�w�.����Y����q9��V�����'�2�o����0���C���]ǻN�����9�%�b��`�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y������b�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�@���N����E
��^ �����u��
���f�W���
����_F�� 1��B���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�j�5�������TF��d:��9�������w�l�W������]ǻN�����9�%�b��o�-����Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�E��e�w�_�u�w�4����	�ѓ�l^��G1�����
�<�u�u���8���B�����Y������m�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�N����l��D��Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�j�5���	����	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�u�W�W���������h,��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�b��n�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lQ��h_�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&Ĺ��V��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�
�e�4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�&�֓�C9��S1�����u��
���}�J���^���F��P ��U���
�
�d�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��7��
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u���(�������W9��h��U����
���l�}�Wϭ�����C9��u1�*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u���(�������TF��d:��9�������w�l�W������]ǻN�����9�%�b��f�����Cӵ��l*��~-��0����}�`�1� �)�W���C���V��^�E��e�e�n�u�w�.����Y����q9��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�b��d�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����q9��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����;����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��B���d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�j�5��&����_��E��Oʆ�����m�}�G��Y����Z��[N��B���d�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h,��A���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b��l�(�������]9��PN�&������_�w�}����Ӗ��l$��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�b��l�(���
���5��h"��<������}�b�9� ���Y����F�D�����
�
�
�`�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�N����9��h��*���&�2�o����0���s���@��V��*݊�
�`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�@����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�d�:���	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l+��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L���d�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ށ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��8���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�
9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ߓ�lT��G1�����
�<�u�u���8���B�����Y������g�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�@����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�d�:���	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l+��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L���a�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ہ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��8���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�
9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ߓ�lS��G1�����
�<�u�u���8���B�����Y������`�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�@����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�d�:���	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l+��h�����%�0�u�u���8���Y���A��N�����4�u�
�
����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L���b�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(؁�	����l��PN�&������o�w�m�L���Yӕ��]��G1��8���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�
9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ߓ�l^��G1�����
�<�u�u���8���B�����Y������m�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�@����l��D��Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�d�:���	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
���(�������]9��PN�&������_�w�}����Ӗ��l+��h�����%�0�u�u���8���Y���A��N�����4�u�
�
��m��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�l��d�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y������d�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�N���Hù��l��h���������g�W��B�����Y������d�
�;�$�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hW��*���%�0�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W���������h#��D���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
��l��������V�=��*����u�h�r�p�W�W���������h#��G���
�<�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����~9��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����&ʹ��T��G1�����
�<�u�u���8���B�����Y������d�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&ʹ��U��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�N���H����V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�d�:��&����_��Y1���������W�W���������h#��F���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�d�:��&����Z�=��*����
����u�FϺ�����O��N�����4�u�
�
��i����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�
�c�<�(���&����Z�=��*����n�u�u�$�:����&ʹ��R��G1�����0�u�u����>���D����l�N�����u�
�
�
�b�4�(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������d�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L���d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�d�:��&����_��E��Oʆ�����m�}�G��Y����Z��[N��*���
�1�
�e�w�}�8���8��ƹF��^	��ʳ�
�!��'��2�(���I����l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l*��G1�*ڊ�=�
�0�
�b�j�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�e�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������U��]��G��������4���Y����\��XN�N���u�&�2�4�w�
���� ����@9��h_�F���u�u��
���(���-���S��X����n�u�u�&�0�<�W�������|��D1����`�u�u����>���<����N��
�����e�n�u�u�$�:����5����u	��{��*ފ�
�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^"�����'��:�
���(���&����\��c*��:���
�����}�������9F������3�
�!��%�����J�ד�[��B1�CҊ�f�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����\��X��Dي�
�=�
�0��h�E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������,� �
�c�f�;�(��L����	F��s1��2������u�f�}�������9F������<�
����)�Fف�&����S��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GU��D��U����
���l�}�Wϭ�����R��^	�����a�u�u����L���Yӕ��]��P�����g�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��]	��h�����'�2�d�l�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����L����q)��r/�����u�<�;�9�0�-����Jù��\��c*��:���
�����l��������l�N�����u��;�1��8���&¹��T9��Y��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��%�"���6����
9��Q��Gي�g�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����g��C1�*ۊ�0�
�c�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�`�3�:�i�Mύ�=����z%��N�����4�u�%�&�0�?���M����|)��v �U���&�2�4�u��1�(���&����lR��h_�� ��l�
�g�o���;���:����g)��Z�����:�e�n�u�w�.����Y����Z9��E1�����
�
�
�0��k�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������V��c1��M���8�b�o����0���s���@��V�����2�7�1�b�o�g�5���<����F�D�����%�&�2�6�2��#���@����l^�=��*����n�u�u�$�:����	����l��hV�U������n�w�}�����ƭ�l��h�����
�!�e�3�:�d�Mύ�=����z%��N�����4�u�%�&�0�?���K����|)��v �U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�g�u�w��;���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��]�Oʗ����_�w�}����Ӈ��@��T��*���&�d�
�&��o�Mύ�=����z%��N�����4�u�%�&�0�?���A����|)��v �U���&�2�4�u�%��(��&����V��T��!�����
����_�������V�=N��U���;�9�4�,�g�k�E���I����g"��x)��N���u�&�2�4�w�/�(߁�I����\��c*��:���
�����l��������l�N�����u�'�
�
�g�����
���5��h"��<������}�w�2����I��ƹF��^	��ʴ�,�e�c�g�4�l�Mύ�=����z%��N�����4�u�'�
��m�(���Y�Ɵ�w9��p'�����u�<�;�9�6�$�G��K����	F��s1��2������u�d�}�������9F������4�,�e�c�e�,�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^"�����'��:�
��8�(��Y�Ɵ�w9��p'��#����u�a�1� �)�W���s���@��V�����2�6�0�
��.�A������5��h"��<��u�u�&�2�6�}��������l^��T��:����n�u�u�$�:��������U��V�����u��
����2���+������Y��E��u�u�&�2�6�}����&¹��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������`2��C_�����d�u�u����>��Y����Z��[N��*���
�1�
�e�w�}�8���8��ƹF��^	��ʳ�
���,�"��(���A�ޓ�F��d:��9�������w�n�W������]ǻN�����9�3�
���$����&����^��N�&���������W��Y����G	�UךU���<�;�9�3���;�������U��V��D��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���5����G9��h_�� ��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����~3��N!��*���d�3�
�g��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U��^��E��������4���Y����W	��C��\�ߊu�u�<�;�;�)����&����CW�=��*����
����u�W������]ǻN�����9�&�9�!�'����@����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d�1��@܁�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
� �o�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���c�3�
�c��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1��ފ� �m�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��Q��Aي�g�o�����4���:����V��X����n�u�u�&�0�<�W�������U��_��G��������4���Y����\��XN�N���u�&�2�4�w�8�$�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��1�(���A�ѓ� F��d:��9�������w�l�W������]ǻN�����9�:�
�:�3����J����	F��s1��2������u�g�9� ���Y����F�D�����'�6�;�g�1��Fځ�K����g"��x)��*�����}�u�8�3���B�����Y�����0�g�3�
�g��D��*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T�� ��&���
� �l�d�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��ي� �l�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V��[Z�� ��b�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����V
��Q��Aۊ�f�o�����4���:����W��S�����|�_�u�u�>�3�ϰ�����l ��[�����u��
����2���+������Y��E��u�u�&�2�6�}����˹��l_��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*��������
9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��1�G���&����CU�=��*����
����u�BϺ�����O��N�����4�u�0��;�l����A¹��\��c*��:���
�����h��������l�N�����u�0��9�e�;�(��&���5��h"��<������}�b�9� ���Y����F�D�����0�
�8�`�1��G���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʦ�9�!�%�
�"�l�Fށ�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�l�3��m�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����!�%�e�3��m�B���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����!�%�d�3��m�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����!�%�g�3��m�N���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����0�c�3�
�c��D��*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T�� ��&���f�3�
�l��n�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��R����
� �d�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�e�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��D݊� �d�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��C���
�e�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_�����e�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��]�� ��c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������R��B1�E݊�f�o�����4���:����W��S�����|�_�u�u�>�3�ϰ�����9��h_�L���u�u��
���(���-���S��X����n�u�u�&�0�<�W�������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}�����ғ�F9��Y��G��������4���Y����\��XN�N���u�&�2�4�w�8�$���O����W��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*���&����R��G]��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u�%�>��������Q��N�&���������W������\F��d��Uʦ�2�4�u�0��1�O���&����l��N��1��������}�F�������V�=N��U���;�9�;�"�2�l�(���H����CU�=��*����
����u�BϺ�����O��N�����4�u�0��;�l����H�ߓ� F��d:��9�������w�l�W������]ǻN�����9�;�"�0�e����Aƹ��\��c*��:���
�����h��������l�N�����u�0��9�d�;�(��H����	F��s1��2������u�f�}�������9F������;�"�0�g��(�F��&���5��h"��<������}�b�9� ���Y����F�D�����0��9�`�1��E���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʻ�"�0�g�
�"�l�Fށ�J����g"��x)��*�����}�`�3�*����P���F��P ��U���
�8�g�
�"�l�E؁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�"�l�D܁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�"�l�C߁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�"�l�C؁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�"�l�Bہ�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�"�l�Aށ�J����g"��x)��*�����}�d�3�*����P���F��P ��U����9�e�3��l�F���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����0�g�
� �f�l�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V����� �m�b�6�w�}�#���6����9F������2�%�3�
�d����*����|!��d��Uʦ�2�4�u�%������Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��*���
�1�
�e�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��d�MϜ�6����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w�-��������Q�,��9���n�u�u�&�0�<�W���
����W��X��U�����n�u�w�.����Y����Z��S
��B���u����l�}�Wϭ�����R��^	�����m�u�u����L���Yӕ��]��V�����1�
�m�o���2���s���@��V�����2�7�1�c�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��k�MϜ�6����l�N�����u�%�&�2�5�9�O���Y����v'��=N��U���;�9�4�
�>�����M����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:����	����l��h_�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�g�u�u���6��Y����Z��[N��*���
�1�
�d�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&���� S��N��:����_�u�u�>�3�Ͽ�&����Q��X�Oʗ����_�w�}����Ӈ��@��U
��G��o�����W�W���������D�����g�f�o����9�ԜY�ƿ�T�������7�1�g�g�m��8���7���F��P ��U���&�2�7�1�e�l�MϜ�6����l�N�����u�%�&�2�5�9�E��CӤ��#��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-��������^�,��9���n�u�u�&�0�<�W���
����W��Y��U�����n�u�w�.����Y����Z��S
��E���u����l�}�Wϭ�����R��^	�����c�u�u����L���Yӕ��]��V�����1�
�`�u�w��;���B�����Y�����<�
�1�
�a�}�W���5����9F������4�
�<�
�3��@���Y����v'��=N��U���;�9�4�
�>�����A����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�M������]�}�W�������C9��P1����b�o�����}���Y����R
��G1�����1�f�c�o���2���s���@��V�����2�7�1�a�b�g�5���<����F�D�����%�&�2�7�3�i�C��;����r(��N�����4�u�%�&�0�?���J����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lR��T��:����n�u�u�$�:����	����l��hZ�U������n�]�}�W���	����GF��r_�1���
�
�8�9�d�3�(���
����9��O1��ʜ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�f�
�3���Cӯ��v!��d��U���u�1� �
��	�W���7����aF�=N��U���!�}�u�u�w�}����Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W�������f2��c*��:���
�����l��������O��N�����6�8�:�0�#�W�}���Y����\��CN��0���e�
�
�>�2���
����F��=N��U���0�<�u�_�w�}�W���=����}2��r<�U���u�u�����2��0����v4��N��U���1�;�
���}�W���<����9F�N��U���!����m��#���+����F�G��U�ߊu�u�u�u�;�}�W���*����|!��d��U���u�'�&�!�m��W���&����p]ǻN��U���<�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������z(��c*��:���n�u�u�u�w�9����Y����`2��{!��6�����u�f�w�2����I���9F���U���%�;�;�n�]�}�WϽ�����]��+�B��3�e�4�,�g�k�Eϗ�s���T��E��]���u�u�u��#�
����Cӯ��v!��d��U���u��1�0�$�<����Y����t#��=N��U���u�1�'�&� �9���0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�1�%�.�G��0�Ɵ�w9��p'��#����u�f�1� �)�W���s���F�T�Oʜ�u��
���f�W���Y����F��x;��&���������W��Y����G	�UךU���u�u�1�'�$�l�Mϗ�Y����)��t1��6���u�f�1�"�#�}�^�ԜY���F��N�<����
���l�}�W���Yӑ��\��yN��1�����_�u�w�}�W��Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N��D��������4���:����U��S�����|�|�_�u�w�3�W���	����G]Ǒ=d�����u�u�4�,�g�k�E���CӅ��C	��Y��@��b�d�3�e�6�$�G��K�����R��U���u�_�u�u�w�}��������X�BךU���u�u�1�'�$�����D����l�N��Uʔ�1�0�&�<�#�}�I��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����E��E��u�'�
�
�g�����
����F�N����h�u�'�
��m�(���U���F��H���'�
�
�e��m�}���Y���R��R��U��4�,�e�c�e�<����
��ƹF�N�����k�4�,�e�a�o���s���F�@�H���'�
�
�e��8�[���Y�����
P�����
�e�
�d�]�}�W���Y���F��N1��C���$�|�_�u�w�;�G�������]�� ��F؊�
�4�
�&��m�MϽ�����]��+�B��3�e�3� ��o�������lW��V���ߊu�u�0�0�>�}����s���F�~*��K��_�u�u�u�w��(���>���W�N��U���1�;�
���}�I��U���F�
��D�����h�u�e�W�W���Y�ƨ�F��~*��U��f�|�u�u�'�/�W���Y���F�N�����k�3�
���$����&����^��BךU���u�u�<�d�j�}�$���,����F��h��M���%�y�u�u�w�}����Y����`9��b"��:���&�3�
�d��o�L�ԜY�ƪ�9��B��G���f�;�
�g�f�0����	����	F��Z�����8��l��g��(�������@9��Y��G���8�-�1�%�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�o�}���Y������FךU���u�u�<�e�j�}�$���,����F��1�����g�
�e�_�w�}�W������F��h��9��� �
�l�d�1��E܁�H���F�N�� ���k�3�
���$����@�ד�F9��1��\�ߠu�u�3�e�$�)����K����lT��N����:�0�!�8��d�3���&ù��G	��h]��*���g�u�u�2�9�/�ϳ�	��ƹF�N��1��u�y�u�u�w�}�9���*����[�BךU���u�u�<�e� ��?��Y����F�N�����
���u�i�n�^���YӖ��GF��GN��U���u�u�6�>�j�}�������F�N�����h�u�%�'�#�W�W���Y�ƨ�]V�	N�����
�g�
�e�]�}�W���Y���F��G1��*��
�0�_�u�w�}�W������T��Q��G݊�d�n�_�u�w��(���������1�� ���u�:�%�;�9�}�B��N����lV��^����&�f�
�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��^ �H���'�
� �m�g�-�[���Y�����
P����� �m�e�6�{�}�W���Yӂ��GF�	��*���m�e�%�|�]�W�}���Y���G��T�����&�4�0�}�'��(���PӉ��G��D��ʸ�6�<�0�u�z�}�WϿ�&����@��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���%��
�&�w�`����-����l ��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�$�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�e��"��m��������V��D��ʥ�:�0�&�u�z�}�WϮ�I����r/��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����z9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�e��"��m��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l4��v'��*���#�1�%�0�w�`����+����lV��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��D'��1�����&�<�;�%�8�8����T�����h<��4���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�I����r/��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�'�m�%���0�֓�C9��SG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P�����YNךU���u�u�u�u�w�}�W���&ù��D'��1�����h�%�e�� ��G�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6��(�������W9��R	�����;�%�:�0�$�}�Z���YӖ��l4��v'��E���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l4��v'��E���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N��U���u�u�u�%�g�� ���Hù��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*����
�e�4��1�(������C9��e��<��
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��'����d�
�'�0�<����Y����V��C�U���%�e��"��l�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*����
�e�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����z9��h�����|�u�=�;�]�}�W���Y���F�N������"��d��/���Y����a��~1�N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��@/��Dۊ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�4���F���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4���F���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$���������� O�C��U���u�u�u�u�w�}�W���Y�����h<��4���d�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�c�t����Y���F�N��U���u�u�u�u�w��(���8����l��A�����u�h�%�e��*�>��&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�%���0����C�������%�:�0�&�w�p�W���	�֓�R��h_�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���8����l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������"��d��-����P�Ƹ�V�N��U���u�u�u�u�w�}����+����lW��G��U��%�e��"��l�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�� ��F݁�	����l��PN�����u�'�6�&�y�p�}���Y����a��~1�*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����a��~1�*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��Dފ�&�
�f�|�#�8�W���Y���F�N��U���u�u�u�
��<�6���K����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9�� G�����_�u�u�u�w�}�W���Y���F�G1��'����d�
�%�!�9����Y����lV��V��*���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h^�����
�g�%�0�w�.����	����@�CךU���
�
�4���o����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��'����d�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����+����lW��V�����|�!�0�u�w�}�W���Y���F�N��*ڊ�4��
�g�'�8�W��	�֓�R��h_����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l4��v'��F���
�9�
�'�0�<����Y����V��C�U���%�e��"��l�(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e��"��l�(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Fہ�
����O��_�����u�u�u�u�w�}�W���Y���C9��e��<��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�d�a�}����s���F�N��U���u�u�u�u�'�m�%���0����R��[
�����i�u�
�
�6��(�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u������&�Փ�A��V�����'�6�&�{�z�W�W���&ù��D'��]�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�m�%���0����C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ڊ�4��
�f�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(߁�����U��E��I���
�
�4���n�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�4���C���&����C�������%�:�0�&�w�p�W���	�֓�R��h_�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�R��h_�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��A���8�d�|�u�?�3�}���Y���F�N��U���u�u�%�e��*�>��&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lW��N�����u�u�u�u�w�}�W���Y���F��h^�����
�a�4�
�;�����E�Ƽ�9��@/��Dފ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����d�
�'�2�6�.��������@H�d��Uʥ�e��"��f���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^�����
�a�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(߁�����R��G1�����u�=�;�_�w�}�W���Y���F�N��E���"��d�
�%�:�K���&ù��D'��Z�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����a��~1�*���#�1�%�0�w�.����	����@�CךU���
�
�4���h��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�4���h��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�w�}�W���Y����lV��V��*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�m�~�)����Y���F�N��U���u�u�u�u������&�ӓ�C9��S1�����h�%�e�� ��Fځ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g�� ���Hƹ��V��D��ʥ�:�0�&�u�z�}�WϮ�I����r/��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&�ӓ�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��E���"��d�
�'�+����Y����l�N��U���u�u�u�u�w�-�G�������9��R	��Hʥ�e��"��f�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�e��"��l��������V��D��ʥ�:�0�&�u�z�}�WϮ�I����r/��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����z9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N��U���%�e��"��l��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l4��v'��*���#�1�%�0�w�`����+����lW��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��D'��1�����&�<�;�%�8�8����T�����h<��4���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�I����r/��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e��"��l���������YNךU���u�u�u�u�w�}�W���&ù��D'��1�����h�%�e�� ��F�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6��(݁�	����l��PN�����u�'�6�&�y�p�}���Y����a��~1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�R��h\�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
�6��(݁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������O��_�����u�u�u�u�w�}�W���Y���C9��e��<���4�
�9�
�%�:�K���&ù��D'��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l4��v'��*���2�4�&�2�w�/����W���F�G1��'����g�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����a��~1�����u�h�4�
�8�.�(���O����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�6��(݁�	����O�C��U���u�u�u�u�w�}�W���YӖ��l4��v'��*���2�i�u�
��<�6���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g�� ���J����E
��G��U���<�;�%�:�2�.�W��Y����lV��V��*ي�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��@/��F���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N��U���u�u�u�%�g�� ���J����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��N�����u�u�u�u�w�}�W���Y���F��h^�����
�
�%�#�3�-����DӖ��l4��v'��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��e��<���%�0�u�&�>�3�������KǻN��*ڊ�4��
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��V��*ي�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�g�� ���J����E
��G�����_�u�u�u�w�}�W���Y���C9��e��<���%�0�u�h�'�m�%���0����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���8����R��[
�����4�&�2�u�%�>���T���F��1�����a�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h<��4���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���u�u�u�u�w��(���8����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hV�U���;�_�u�u�w�}�W���Y���F�N��E���"��a�4��1�(������C9��e��<���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h^�����
�
�'�2�6�.��������@H�d��Uʥ�e��"��c�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����a�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(���8����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h^�����
�
�'�2�k�}�(߁�����]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����+����lS��G1�����0�u�&�<�9�-����
���9F���*����
�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��'����`�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�l�^������F�N��U���u�u�u�u�w�}����+����lS��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��L���!�0�u�u�w�}�W���Y���F�N��U���
�4��
��-����	����[��h^�����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���"��`�%�2�}����Ӗ��P��N����u�
�
�4���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*����
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����+����lS��G1�����u�=�;�_�w�}�W���Y���F�N��E���"��`�%�2�}�JϮ�I����r/��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��D'��1��*���
�'�2�4�$�:�W�������K��N������"��c�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�4��
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ù��D'��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����e�|�!�0�w�}�W���Y���F�N��U���u�
�
�4���(�������A��S��*ڊ�4��
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e��"��a�-����
������T��[���_�u�u�
��<�6���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4��
��/���Y����\��h��C��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�֓�R��hX�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e��"��a�-����DӖ��l4��v'��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��@/��B���
�9�
�'�0�<����Y����V��C�U���%�e��"��j��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�4�����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��@/��B���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�d�|�#�8�W���Y���F�N��U���u�u�u�
��<�6���&����_��E��I���
�
�4����������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�� ��@����ƭ�@�������{�x�_�u�w��(���8����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�4���(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��V��*݊�%�#�1�|�w�5��ԜY���F�N��U���u�%�e�� ��@��������h<��4���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����m�4�
�9��/�Ͽ�
����C��R��U���u�u�%�e��*�>�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�6��(ׁ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����U����ߊu�u�u�u�w�}�W���Y���F��1�����m�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�e�t����Y���F�N��U���u�u�u�u�w��(���8����R��[
�����i�u�
�
�6��(ׁ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g�� ���A����TF��D��U���6�&�{�x�]�}�W���&����z9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��<�6���&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h^�����
�
�%�#�3�t�W������F�N��U���u�u�u�%�g�� ���A����TF���*����
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���"��l�4��1�(���Ӈ��Z��G�����u�x�u�u�'�m�%���0�ߓ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u������&ʹ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��]��U���;�_�u�u�w�}�W���Y���F�N��E���"��l�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��D�������9F�N��U���u�u�u�u�w�}�W���&����z9��V�����'�2�i�u������&ʹ��l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�G�������l��PN�����u�'�6�&�y�p�}���Y����a��~1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���8����C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ڊ�4��
�
�'�+����Y����l�N��U���u�u�u�u�w�-�G�������l��PN�U���
�4��
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b��e�4��1�(���Ӈ��Z��G�����u�x�u�u�'�j�5�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�l�(���&�����YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����g�|�!�0�w�}�W���Y���F�N��U���u�
�
�
��-����	����[��hY��*ڊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��E���0�u�&�<�9�-����
���9F���*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N����l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������e�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u���(߁����F�� 1��E�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��h_�����9�
�'�2�6�.��������@H�d��Uʥ�b��d�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&�֓�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��_�U���;�_�u�u�w�}�W���Y���F�N��B���d�
�%�#�3�-����DӖ��l$��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l$��1�����&�<�;�%�8�8����T�����h,��E���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�&�֓�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���d�
�%�#�3�t�W������F�N��U���u�u�u�%�`��F߁����F�� 1��D��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��u1�*���#�1�%�0�w�.����	����@�CךU���
�
�
�d�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�a�3�:�l�^������F�N��U���u�u�u�u�w�}����;����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h]�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�
�d�4�
�;�����E�Ƽ�9��_�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��_�����4�&�2�u�%�>���T���F�� 1��Dۊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����;����C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*݊�
�d�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u���(���	����[��hY��*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h,��G���
�9�
�'�0�<����Y����V��C�U���%�b��d��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������d�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��D�������9F�N��U���u�u�u�u�w�}�W���&����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�F���=�;�_�u�w�}�W���Y���F�N������d�
�%�!�9����Y����lQ��h_�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��h_�����u�&�<�;�'�2����Y��ƹF��hY��*���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������d�
�%�!�9�^������F�N��U���u�u�u�u�'�j�5��&����Z�G1��7��n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��Dي�%�#�1�%�2�}����Ӗ��P��N����u�
�
�
�d�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�f�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�a�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�N���� 9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��A���!�0�u�u�w�}�W���Y���F�N��U���
�
�f�4��1�(������C9��u1�*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��u1�*���2�4�&�2�w�/����W���F�G1��7��
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N���� 9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�f�4��1�^�������9F�N��U���u�u�u�u�w��(���J����TF���*���f�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hY��*���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�b��f���������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��d�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��R��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��F��u�=�;�_�w�}�W���Y���F�N��Uʥ�b��d�
�'�+���������h,��A���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h,��A���0�u�&�<�9�-����
���9F���*���a�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��R��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�b��d�
�'�+����Y����l�N��U���u�u�u�u�w�-�@���Hǹ��V�
N��B���d�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��7��
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
��h��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�`�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�c�;���P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�`�6��������F�� 1��Dߊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��Dߊ�'�2�4�&�0�}����
���l�N��B���d�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�lW��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�`�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(؁�&�ӓ�A��S��*݊�
�`�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��d�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�a�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�N����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�A���=�;�_�u�w�}�W���Y���F�N������d�4�
�;�����E�Ƽ�9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l$��h��ʴ�&�2�u�'�4�.�Y��s���C9��u1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*ۊ�%�#�1�|�w�5��ԜY���F�N��U���u�%�b��f�-����DӖ��l$��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��9��h��*���2�4�&�2�w�/����W���F�G1��7���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��h\�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����K���G��d��U���u�u�u�u�w�}�W���YӖ��l$��h�����%�0�u�h�'�j�5�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(݁�����@��YN�����&�u�x�u�w�-�@���K����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��g�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hY��*؊�'�2�i�u���(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��n��������V��D��ʥ�:�0�&�u�z�}�WϮ�N����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����_�u�u�u�w�}�W���Y���F�G1��7���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�`�~�)����Y���F�N��U���u�u�u�u���(܁�	����l��PN�U���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����f�%�0�w�.����	����@�CךU���
�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��h]�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b��d�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����C��R������f�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��a�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�a�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�N����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�D���=�;�_�u�w�}�W���Y���F�N������a�4�
�;�����E�Ƽ�9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l$��h��ʴ�&�2�u�'�4�.�Y��s���C9��u1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*ފ�%�#�1�|�w�5��ԜY���F�N��U���u�%�b��c�-����DӖ��l$��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��9��h��*���2�4�&�2�w�/����W���F�G1��7���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��h[�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����K���G��d��U���u�u�u�u�w�}�W���YӖ��l$��h�����%�0�u�h�'�j�5�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(ځ�����@��YN�����&�u�x�u�w�-�@���L����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��`�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hY��*ߊ�'�2�i�u���(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��k��������V��D��ʥ�:�0�&�u�z�}�WϮ�N����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����_�u�u�u�w�}�W���Y���F�G1��7���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�b�~�)����Y���F�N��U���u�u�u�u���(ف�	����l��PN�U���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����c�%�0�w�.����	����@�CךU���
�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��hX�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b��a�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����C��R������c�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��b�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�a�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�N����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�M���=�;�_�u�w�}�W���Y���F�N������b�4�
�;�����E�Ƽ�9�� 1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l$��h��ʴ�&�2�u�'�4�.�Y��s���C9��u1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*݊�%�#�1�|�w�5��ԜY���F�N��U���u�%�b��`�-����DӖ��l$��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��9��h��*���2�4�&�2�w�/����W���F�G1��7���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��hV�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����K���G��d��U���u�u�u�u�w�}�W���YӖ��l$��h�����%�0�u�h�'�j�5�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(ׁ�����@��YN�����&�u�x�u�w�-�@���A����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��m�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hY��*Ҋ�'�2�i�u���(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��d��������V��D��ʥ�:�0�&�u�z�}�WϮ�N����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����_�u�u�u�w�}�W���Y���F�G1��7���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�e�~�)����Y���F�N��U���u�u�u�u���(ց�	����l��PN�U���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����l�%�0�w�.����	����@�CךU���
�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��hW�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b��n�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����C��R������l�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�l��e�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�a�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�@����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�L���=�;�_�u�w�}�W���Y���F�N������e�4�
�;�����E�Ƽ�
9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��h��ʴ�&�2�u�'�4�.�Y��s���C9��z1�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hW��*ڊ�%�#�1�|�w�5��ԜY���F�N��U���u�%�l��g�-����DӖ��l+��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ʹ��V��G1�����0�u�&�<�9�-����
���9F���*���e�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#��E���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N��U���u�u�u�%�n��F߁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������_�C��U���u�u�u�u�w�}�W���Y�����h#��E���
�9�
�'�0�a�W���&����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����l��PN�����u�'�6�&�y�p�}���Y����~9��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�n��F߁����F��h�����#�g�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h#��E���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�
�g�-����DӖ��l+��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�lW��V�����'�2�4�&�0�}����
���l�N��L���d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1��Dۊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�f�~�)����Y���F�N��U���u�u�u�u���(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����P�����ߊu�u�u�u�w�}�W���Y���F��1��Dۊ�%�#�1�%�2�}�JϮ�@����9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�@����9��R	�����;�%�:�0�$�}�Z���YӖ��l+��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(���	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��Dۊ�%�#�1�|�w�5��ԜY���F�N��U���u�%�l��f�����E�Ƽ�
9��_�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����~9��h�����%�0�u�&�>�3�������KǻN��*ӊ�
�g�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hW��*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���a�3�8�d�~�}����s���F�N��U���u�u�u�u�'�d�:��&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR��N�����u�u�u�u�w�}�W���Y���F��hW��*���4�
�9�
�%�:�K���&ʹ��T��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ʹ��T��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��\�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�d�:��&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hW��*���4�
�9�|�~�)����Y���F�N��U���u�u�
�
��o����Y����l_��h_����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��1��*���
�'�2�4�$�:�W�������K��N������d�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��8��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���u�u�u�u�w��(���J����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��8��
�%�#�1�'�8�W��	�ߓ�lW��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�lW��G��U���<�;�%�:�2�.�W��Y����l_��h_�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���J����TF������!�9�f�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��8��
�%�#�1�~�}����s���F�N��U���u�u�%�l��l�(������C9��z1�N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��Z�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�
�a�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���a�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�a�3�8�f�t�W������F�N��U���u�u�u�u�w�-�N���Hǹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��[�����u�u�u�u�w�}�W���Y���F���*���a�4�
�9��/���Y����~9��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����~9��h��ʴ�&�2�u�'�4�.�Y��s���C9��z1�*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�N���Hǹ��V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���a�4�
�9�~�t����Y���F�N��U���u�u�u�
���C��������h#��A�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����l_��h_�����9�
�'�2�6�.��������@H�d��Uʥ�l��d�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��L���d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ց�&�ӓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���Y���F�N��L���d�
�%�#�3�-����DӖ��l+��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��1�����&�<�;�%�8�8����T�����h#��@���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ց�&�ӓ�A��S�����;�!�9�f��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��L���d�
�%�#�3�t�W������F�N��U���u�u�u�%�n��Fځ����F��1��D��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��z1�����9�
�'�2�6�.��������@H�d��Uʥ�l��d�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lU��N�����u�u�u�u�w�}�W���Y���F��hW��*ۊ�%�#�1�%�2�}�JϮ�@����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����C�������%�:�0�&�w�p�W���	�ߓ�lW��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��l����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�
9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�
�'�0�a�W���&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�N���K����E
��G��U���<�;�%�:�2�.�W��Y����l_��h\�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y���F�N��Uʥ�l��g�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��O�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�
�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l��e�-����
������T��[���_�u�u�
���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��1�����h�%�l��e�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��n��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�w�}�W���Y����l_��h]�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����f�c�u�=�9�W�W���Y���F�N��U���u�%�l��d�<�(���&����Z�G1��8���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hW��*ي�'�2�4�&�0�}����
���l�N��L���f�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ�� 9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�d�:���	����[��hW��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��z1�����9�
�'�2�6�.��������@H�d��Uʥ�l��a�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR��N�����u�u�u�u�w�}�W���Y���F��hW��*ފ�%�#�1�%�2�}�JϮ�@����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����C�������%�:�0�&�w�p�W���	�ߓ�lR��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��i����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�
9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�
�'�0�a�W���&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�N���L����E
��G��U���<�;�%�:�2�.�W��Y����l_��h[�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y���F�N��Uʥ�l��`�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��F�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�
�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l��b�-����
������T��[���_�u�u�
���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��1�����h�%�l��b�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��k��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�w�}�W���Y����l_��hX�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����a�f�u�=�9�W�W���Y���F�N��U���u�%�l��a�<�(���&����Z�G1��8���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hW��*܊�'�2�4�&�0�}����
���l�N��L���c�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�d�:���	����[��hW��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��z1�����9�
�'�2�6�.��������@H�d��Uʥ�l��b�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�d�t����Y���F�N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR��N�����u�u�u�u�w�}�W���Y���F��hW��*݊�%�#�1�%�2�}�JϮ�@����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����C�������%�:�0�&�w�p�W���	�ߓ�lQ��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��j����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�
9�� 1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�
�'�0�a�W���&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�N���A����E
��G��U���<�;�%�:�2�.�W��Y����l_��hV�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�=�;�_�w�}�W���Y���F�N��Uʥ�l��m�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��C�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�
�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l��o�-����
������T��[���_�u�u�
���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��1�����h�%�l��o�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��d��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�w�}�W���Y����l_��hW�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����a�e�u�=�9�W�W���Y���F�N��U���u�%�l��n�<�(���&����Z�G1��8���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hW��*ӊ�'�2�4�&�0�}����
���l�N��L���l�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��
9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�
�%�!�9�^������F�N��U���u�u�u�u�'�d�:���	����[��hW��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���Z*��^1�����:�
�
�0��m�W�������A	��D�X�ߊu�u��9��2�(���	�ғ�V��[�����;�%�:�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���R��^	�����e�|�!�0�w�}�W���Y���F�N��U���9�
�:�
�8�-�C�������Z�V�����
�#�
�n�w�}�W���Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�c�3�8�b�t����Y���F�N��U���u�u�u��;���������l��hV�U��<�
�<��%�����&¹��A��X�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�;�u�3�w�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����P	��1��*��
�g�h�4��2����¹��O��_��U���u�u�u�u�w�}��������l*��G1�*ڊ�=�
�0�
�b�j�K���*����u	��{��*���e�%�<�3��m�A���B���F�N��U���u��9�
�8�����H����C��E��D��u�h�3�
�#���������lW��_�� ��c�
�f�_�w�}�W���Y���F��h��3����:�
�
������L���F������:�
�:�%�c�l����&����l��G�U���<�
�<��%�����&¹��A��[�]���i�u��9��2�(���	�ғ�l��B1�@ӊ�g�g�n�u�w�4�(���?����\	��1�����2�d�`�}�~�a�W�������A9��X��*ۊ�
� �d�`��o�D��Y���F�N��U����-� �,�"��A�������P��S��"��� �,� �
�a�l����K�ӓ�]ǻN��U���u�u�u�u� �%�"�������A��[�U��<�
����)����&����l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�a�1�0�D���Y����9F�N��U���u�u�u��9�9�(�������9��P1�L���h�2�%�3��n�(��s���F�N��U���3�
�:�0�#�/�(�������
T�
N�����
�g�
�d�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GS��D��\���!�0�_�u�w�}�W���Y���U5��z;�����
�l�d�'�0�l�G���DӀ��K+��c����
�
� �m�d�-�L���Y���F�N��U���9�
�:�
�8�-�C���H����lW�� N�U���9�
�:�
�8�-�C���H����T��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���Z*��^1�����:�
�
�
��8�(��N���[�I����u�x�!�0�9�%�W�������C9��h��\ʺ�u�=�u�!�#�}�������l�N��*���3�8�4�&�0�����CӖ��P��F��*���3�8�u�%�4�q��������W9��B�����:�1�
� �o�n����Y����V��=N��U���u�4�0�4���������F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���
����W��X��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���u�u�9�0�w�}�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�u�u�2�9���Y���F�N�����4�
��&�e�;���D��ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������U��]��G��4�
�:�&��+�(���P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�f�3�:�o�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��F���8�g�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�C�������F�N��U���"�0�u�%���ہ�
����X�N��U���u�u�u�u�6��$������R��c1��@���8�a�_�u�w�}�W���Y������d:��ߊ�&�
�u�k�]�}�W���Y���F�V��&���8�i�u�%���ف�
����9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�-�9���
�����d:��؊�&�
�n�u�w�}�W���Yӑ��]F��h=�����3�8�c�h�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�<�(������F��h=�����3�8�m�_�w�}�W���Y�ƻ�V��G1��*���
�&�
�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���I����l_��N��U���u�u�"�0�w�-�$����֓�@��S����u�u�u�u�w�}�W���7����^F���&���!�d�3�8�f�f�W���Y���F��_������&�d�
�$��G��Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}� ���Y����g9��\�����d�h�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�<�(������F��h=����
�&�
�f�]�}�W���Y���D����&���!�a�3�8�f�}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�?�3�������FǻN��U���u�u�u�u�'��(���Y���k>��o6��-����w�_�u�w�}�W���Y����l�N��ʥ�:�0�&�_�w�}�Z���	����VF��D��U���6�&�{�x�]�}�W�������R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�a�3�8�f�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��D���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���<�9�u�&�>�3�������KǻN�����9�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Qۈ��N��h�����:�<�
�u�w�-��������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W�������[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��S�����;�%�:�0�$�}�Z���YӇ��A��N1�����
�'�6�o�'�2��������F��h��*���$��
�!�c�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���F��R ��U���u�u�u�u�6�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�0�1�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����V��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����a��~1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�f�n�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ڊ�4��
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����W��V�����'�6�&�{�z�W�W���	����l��h_�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h<��4���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e��"��j�������9F���U���6�&�n�_�w�}�Z���	����l��h_�U���<�;�%�:�2�.�W��Y����C9��P1����d�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��E���"��m�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��<�6���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����e�4�&�2�w�/����W���F�V�����1�
�f�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4����������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�G�������l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�f�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�d��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e��*�>��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�֓�R��h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�l�OϿ�
����C��R��U���u�u�4�
�>�����M˹��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(߁�����W��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�a�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����d�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l4��v'��G���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�@��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�4��
�e�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��X�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��'����d�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�e��*�>��&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����`�4�&�2�w�/����W���F�V�����1�
�b�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�4���i������ƹF��R	�����u�u�u�u�w�}�W���
����W�� [��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(߁�����R��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�m�w�.����	����@�CךU���%�&�2�7�3�l�C���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�g�� ���Hƹ��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����a�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l4��v'��@���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����g�`�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��h^�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��n�W�������A	��D�X�ߊu�u�%�&�0�?���M����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@���H����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����q9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�d�<����Y����V��C�U���4�
�<�
�3��C܁�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(݁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�F��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�`�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�o��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�b��n������ƹF��R	�����u�u�u�u�w�}�W���
����W��\��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�&����l��G�U���0�1�%�:�2�.�}�ԜY�����D�����g�d�4�&�0�}����
���l�N��*���
�1�
�c��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����P��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�5�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�g�e�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b��`�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Lʴ�&�2�u�'�4�.�Y��s���R��^	�����b�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*݊�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����N���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b��a�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��V�����;�%�:�0�$�}�Z���YӇ��@��U
��G���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��7���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�E��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����_��V�����'�6�&�{�z�W�W���	����l��h\�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h,��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��d�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������m�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������lU��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��F���h�}�%���.�_�������V�
N��*���&�
�#�
�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����I�ƭ�@�������{�x�_�u�w�-��������P��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ѓ�l_��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�e�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F�� 1��L���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�D������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�d�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��u1�*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��E���
������T��[���_�u�u�%�$�:����J�ғ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����;����R��[
��U���7�2�;�u�w�}�W���Y�����D�����f�a�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�DϿ�
����C��R��U���u�u�4�
�>�����J����@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(؁�&�ԓ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����f�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��\�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��i�W�������A	��D�X�ߊu�u�%�&�0�?���K����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@���H����l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����g�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l$��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�d�l�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(���M����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����q9��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�a�}����Ӗ��P��N����u�%�&�2�5�9�D�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�j�5��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��F��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ѓ�lW��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�f�n�<����Y����V��C�U���4�
�<�
�3��Aց�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(߁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�@����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�b�u�$�4�Ϯ�����F�=N��U���&�2�7�1�d�e��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�l��l������ƹF��R	�����u�u�u�u�w�}�W���
����W�� V��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�&¹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����f�b�4�&�0�}����
���l�N��*���
�1�
�m��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&���� ^��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�c�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�l��f�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�@ʴ�&�2�u�'�4�.�Y��s���R��^	�����e�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ӊ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����I���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�l��c�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Z�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��8���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�C��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����T��V�����'�6�&�{�z�W�W���	����l��hZ�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h#��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��o�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������c�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�
9�� 1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�e�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������W��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ߓ�l^��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�a�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��M���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����a�e�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����l_��hW�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��h�W�������A	��D�X�ߊu�u�%�&�0�?���@����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�N���Hù��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����l�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l+��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�c�e�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(���H����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����~9��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�`�}����Ӗ��P��N����u�%�&�2�5�9�C�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�d�:��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��A��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ�lW��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�a�a�<����Y����V��C�U���4�
�<�
�3��Oف�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��M���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ʹ��U��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�l�6�.��������@H�d��Uʴ�
�<�
�1��d��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e��*�>�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��L��u�}�%�6�9�)���������h<��4���
�%�#�1�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�n�}����Ӗ��P��N����u�%�&�2�5�9�C�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�d�:��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��A���i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ�lW��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�`�c�<����Y����V��C�U���4�
�<�
�3��Gہ�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��E���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ʹ��S��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�m�6�.��������@H�d��Uʴ�
�<�
�1��e��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e��*�>�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��M��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�I����r/��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�g�}����Ӗ��P��N����u�%�&�2�5�9�A�������]9��X��U���6�&�}�%�$�<����&ù��D'��1��*���
�;�&�2�w��(���8����R��[
�����2�u�
�
�6��(݁�	����l��D��U���
�4��
��-��������TJ��h^�����
�
�%�#�3�4�(���UӖ��l4��v'��*���#�1�<�
�>�q����+����lP��G1�����
�<�y�%�g�� ���N����E
��^ �����%�e��"��e��������l��N��E���"��l�4��1�(���
���C9��e��<��
�%�#�1�>����	�֓�R��h_�����9�
�;�&�0�}�(߁�����T��G1�����
�<�y�%�g�� ���H����l��h�����u�
�
�4���C���&����Z��^	�����"��d��-��������TJ��hY��*ڊ�%�#�1�<��4�[Ϯ�N����l��A�����<�y�%�b��o��������l��N��B���f�4�
�9��3����Y����q9��V�����;�&�2�u���(ځ�	����l��D��U���
�
�
�%�!�9��������lQ��hY�����1�<�
�<�{�-�@���A����E
��^ �����%�b��l�6���������F�� 1��Dڊ�%�#�1�<��4�[Ϯ�N����9��h��*���&�2�u�
���E���&����Z��^	�����d�
�%�!�9��������lQ��h_�����9�
�;�&�0�}�(؁�&�ӓ�C9��S1��*���y�%�l��g�<�(���&����Z�G1��8���4�
�9�
�9�.����&ʹ��9��h��*���&�2�u�
���(�������]9��PB��*ӊ�
�
�%�#�3�4�(���UӖ��l+��h�����<�
�<�y�'�d�:�������W9��h��Yʥ�l��b�4��1�(���
���C9��z1�����9�
�;�&�0�}�(ց�&ʹ��l��h�����u�
�
�
�g�<�(���&����Z�G1��8��
�%�#�1�>����	�ߓ�lW��V�����;�&�2�u���(�������W9��h��Yʥ�l��d�
�'�+����&������h#��@���
�9�
�;�$�:�}���Y����]l�N��U���u�u�u�4��4�(���&����[���*���
�%�#�1�>�����Y����\��h�����|�:�u�%�n��F���&����Z��^	��U���6�;�!�9�0�>�G����μ�
9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�
�'�+����&����F��h�����:�<�
�|�8�}����4�ғ�C9��S1��*���u�u�%�6�9�)�������\�G1��8���4�
�9�
�9�.�������]��[����u�'�}�
���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l+��h�����<�
�<�u�w�-��������Z��N��U¥�l��m�4��1�(���
�����T�����2�6�e�u�%�u�(ց�&ʹ��l��h�����h�4�
�:�$�����&����AF��hW��*���4�
�9�
�9�.�������]��[����u�'�}�
���F���&����Z��^	��U���6�;�!�9�0�>�G����μ�
9��\�����1�<�
�<�w�}��������\��h^�����%�l��d��-��������TF�V�����
�:�<�
�~�2�WǮ�@����9��h��*���&�2�h�4��2��������O��EN��*ӊ�
�`�4�
�;���������C9��Y�����6�e�u�'���(���&����_��Y1����4�
�:�&��2����PӉ����h,��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b��e�<�(���&����Z������!�9�2�6�g�}����&Ĺ�� 9��h��*���&�2�h�4��2��������O��EN��*݊�
�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�j�5�������W9��h��U���%�6�;�!�;�:���Y���C9��u1�����9�
�;�&�0�`��������_	��T1�U���}�
�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�N����l��A�����<�u�u�%�4�3��������F��F��B���l�4�
�9��3����DӇ��P	��C1�����e�u�'�}���(�������W9��h��U���%�6�;�!�;�:���Y���C9��u1�*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b��f���������@��
N��*���&�
�:�<��t����	�ѓ�lW��V�����;�&�2�h�6�����&����P9����]���
�
�a�4��1�(���
�����T�����2�6�e�u�%�u�(؁�&�ӓ�C9��S1��*���u�u�%�6�9�)�������\�G1��'����e�4�
�;���������C9��Y�����6�e�u�'���(���8����R��[
�����2�h�4�
�8�.�(�������	����*����
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G�������l��A�����<�u�u�%�4�3��������F��F��E���"��a�4��1�(���
�����T�����2�6�e�u�%�u�(߁�����9��h��*���&�2�h�4��2��������O��EN��*ڊ�4��
�
�'�+����&����F��h�����:�<�
�|�8�}����+����lQ��G1�����
�<�u�u�'�>��������lV�X������"��m�6���������[��G1�����9�2�6�e�w�/�_���&����z9��V�����;�&�2�h�6�����&����P9����]���
�4��
�g�<�(���&����Z������!�9�2�6�g�}����&ù��D'��_�����1�<�
�<�w�}��������\��h^�����%�e��"��l�(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l4��v'��F���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�6��(�������W9��h��U���%�6�;�!�;�:���Y���C9��e��<��
�%�#�1�>�����Y����\��h�����|�:�u�4��)����Y����\��h�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�a�d�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��4�(�������@��Q��E���%�&�2�7�3�k�A�ԜY�Ʈ�T��N��U���u�u�u�u�6���������
F�F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}����	����l��hX�\��u�u�0�1�'�2����s���F������7�1�c�u�$�4�Ϯ�����F�=N��U���&�2�7�1�a���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�6��(݁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����z9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�b�e�<����Y����V��C�U���4�
�<�
�3��F݁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�b�g�<����Y����V��C�U���4�
�<�
�3��C߁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�b�e�<����Y����V��C�U���4�
�<�
�3��B݁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&���� F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�b�w�.����	����@�CךU���%�&�2�7�3�j�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��<�6���&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��B���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ù��D'��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�`�i�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����P��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�`�k�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����Q��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�`�e�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����^��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�m�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����V��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�o�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����W��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�i�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����T��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�e�AϿ�
����C��R��U���u�u�4�
�>�����JŹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��_�����:�d�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�O������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����z9��V�����u�u�7�2�9�}�W���Y���F������7�1�m�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����a�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����A����@��YN�����&�u�x�u�w�<�(���&����Q��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��M��i�u�4�
�8�.�(���&���R��d1�����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����@����@��YN�����&�u�x�u�w�<�(���&����
V��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��L��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������l_��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����a��~1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�n�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��E���"��`�4��1�^��Y����]��E����_�u�u�x�w�-��������`2��C_�����l�4�&�2�w�/����W���F�V�����&�$��
�#�m����@����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:�����3�8�l�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��D���8�d�u�&�>�3�������KǻN�����2�6�0�
��.�Fށ�
����l��^	�����u�u�'�6�$�u��������l^��d��Uʷ�2�;�u�u�w�}��������T9��S1�A���=�;�_�u�w�}�W���Y����Z��D��&���!�d�3�8�f�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�l����H�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�g�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��_�����;�%�:�u�w�/����Q����Z��S
��F���u�u�7�2�9�}�W���Yӏ����D�����m�c�u�=�9�W�W���Y���F��h��*���$��
�!�e�;���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���K����lW��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!�d�;���Y����T��E�����x�_�u�u�'�.��������l��1����
�&�<�;�'�2�W�������@N��h��*���
�a�|�u�w�?����Y���F��QN�����2�7�1�m�o�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����U��D��G��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���������� F��D��U���6�&�{�x�]�}�W���
����@��d:�����3�8�d�
�$�4��������C��R�����<�
�1�
�g�t�W�������9F�N��U���}�%�&�2�5�9�N��Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(���&����l5��D�*���
�f�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����U��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�
�&�
��.����	����	F��X��´�
�<�
�1��m�}���Y����]l�N��Uʼ�u�4�
�<��9�(��Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���&����F��D��U���6�&�{�x�]�}�W���
����@��d:��؊�&�
�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�d�~�}�Wϼ���ƹF�N�����%�&�2�7�3�j�E������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���܁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�a�|�w�}�������F���]���&�2�7�1�`�m�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*���� 9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�(���&�ƭ�@�������{�x�_�u�w�-��������`2��CZ�����
�&�<�;�'�2�W�������@N��h��*���
�`�|�u�w�?����Y���F��QN�����2�7�1�b�e�}����s���F�N�����<�
�&�$���ہ�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*ފ�&�<�;�%�8�}�W�������R��^	�����c�|�u�u�5�:����Y����������7�1�b�a�w�5��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$���ƹ��^9��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����GP��D��*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�m�f�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l ��hX�����;�%�:�u�w�/����Q����Z��S
��B���u�u�7�2�9�}�W���Yӏ����D�����b�c�u�=�9�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$���؁�
����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�
�&��}����Ӗ��P��N����u�%�&�2�4�8�(���
�ޓ�@��h�����%�:�u�u�%�>����	����l��hY�\���u�7�2�;�w�}�W�������C9��P1����m�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���@����l^��D�����:�u�u�'�4�.�_���
����W��^��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��M��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������V��V
�����u�&�<�;�'�2����Y��ƹF��E��*��
�1�'�&�g�<����&����\��E�����%�&�2�6�2��#���K����lW�V�����&�$��
�#�����UӇ��@��T��*���&�m�3�8�`�}��������B9��h��*���
�y�4�
�>�����*����V��D��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�l�(���&���R��^	������
�!�f�1�0�F���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�n����H���G��d��U���u�u�u�4�.�m�A�������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����W����ߊu�u�u�u�w�}����&����R��R��U��4�
�:�&��+�C���M�����Y��E��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������lP��h�����e�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�!�0�u�w�}�W���Y����A��hX�*���'�&�e�i�w�-��������9��N�Dʱ�"�!�u�|�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��N1��C���4�1�0�&�w�`��������_��hX��U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�b�|�#�8�W���Y���F���*ڊ�e�
�1�'�$�m�K���	����@��AX��A��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����e�c�g�4�3�8����DӇ��P	��C1��Cފ�}�u�u�u�8�3���B���F������}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�^Ϫ���ƹF�N��U���'�
�
�e��9����I���R��X ��*���a�e�a�x�f�9� ���Y����F�N�����u�u�u�u�w�}�WϿ� �֓�T��S
����i�u���u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��1�G���1�0�&�u�$�4�Ϯ�����F�=N��U���
�
�e�
�3�/��������]9��X��U���6�&�}�%�$�:����&����GT��D��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�`�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1�U���&�2�6�0��	���&����V�V�����&�$��
�#�o����H����C9��P1������&�d�
�$��E���	����l��F1��*���
�&�
�y�#�-�F���&����l����*܊�
� �d�e��l�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�c�1�0�B�������9F�N��U���u�'�
�
�g�����
���F��G1��D���
�f�e�%��}�W�������V�=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�B��������YNךU���u�u�u�u�%��(��&����V��R�����d�3�
�g�n�-�_���Y�ƨ�D��^����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���H����^9��G�����_�u�u�u�w�}�W���&ù��9��S�����h�4�
�:�$�����?���W��X����n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���!�0�u�u�w�}�W���YӇ��lV��\�����&�d�i�u�'�>��������wN��N����!�u�|�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�=�9�W�W���Y���F��N1��C���4�1�0�&�w�`��������_��h,��U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�w�5��ԜY���F�N�����c�g�4�1�2�.�W������]��[�*���u�u�u�:�9�2�G��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�l�3�8�o�t����Y���F�N��U���
�
�e�
�3�/���E�ƭ�l��D�����b�a�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���4�,�e�c�e�<����
�����T�����c�
�}�u�w�}�������9F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�`�;���PӒ��]FǻN��U���u�u�'�
��m�(�������Z�V�����
�#�a�f�c�p�FϺ�����O��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�4�.�m�A�������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�0�]�}�W���Y���R��1�G���1�0�&�u�j��/���B���F���U���u�u�u�0�3�-����
��ƓF�C�����
�e�
�0�w�.����	����@�CךU���'�
�
�e��8�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����y�4�
�<��.����&����U��B�����2�6�0�
��.�O������R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�y�6�����
����g9��_�����e�u�%�&�0�>����-����9��Z1�Yʴ�
�<�
�&�&��(���J����lW��=N��U���<�_�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�b�3�8�a�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��E���PӒ��]FǻN��U���u�u�'�
��m�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�,�e�c�g�4�m�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<����O�ԓ�VW��D��ʥ�:�0�&�u�z�}�WϿ� �֓�T��R_�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����c�u�%�&�0�>����-����l ��hY����<�
�&�$���ց�
������D�����
��&�d��.�(������T9��R��!���d�
�&�
�g�}��������B9��h��G���8�d�y�4��4�(�������@��h��*��u�%�&�2�4�8�(���
�Г�@��d��Uʷ�2�;�u�u�w�}����Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h_��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�`�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��^��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�g�3�:�l�^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����U��D��G���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�c�1�0�B���PӒ��]FǻN��U���u�u�'�
��m�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�,�e�c�g�4�l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<����O�ԓ�F��D��U���6�&�{�x�]�}�W���&ù��9��h�����%�:�u�u�%�>����*����2��B��L���'�2�d�e�{�<�(���&����l5��D�����a�u�%�&�0�>����-����l ��h[������,� �����A����9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�<����O�ԓ�F��������!�d������O����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�4�,�e�a�o����DӀ��K+��c�����3�
�d�
�e�W�W���Y�Ʃ�@�N��U���u�u�4�,�g�k�E���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�,�e�c�e�*�FϿ�
����C��R��U���u�u�4�,�g�k�E���H����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=�����3�8�a�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C[�����|�u�'�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P���G��d��U���u�u�u�4�.�m�A������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�'�
�
�g�����DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�%����¹��l^��h�I���d�u�=�;����������\��h��*��u�u�%�6�9�)����H����_��^�����u��9�
�8�����H����C��Q��E���%�u�h�_�w�}�W���&ʹ��9��h��U���;�}�0�
�:�n����Nʹ��V�
N��R���9�0�_�u�w�}�W���&����9��h_�L���n�u�u�3��)�1���5����U��h��*���d�c�
�f�k�}�W���Y����l_��h_�����2�"�0�u�$�1����@����W��h�E���u�d�|�0�$�}�W���Y����V
��Z�*���d�c�
�f�]�}�W�������J)��h_��D���
�g�
�e�k�}�$���&����	��h_��D���<�'�2�d�a�f�W�������f*��x��Dӊ�
� �m�f�'�}�Jϸ�&����l��Z1�*ۊ�0�
�`�b�]�}�W�������J)��h�� ��m�%�u�h�1���������C9��h^�����0�
�`�b�]�}�W�������J)��h�� ��m�%�u�h�1���������@9��P1�L��_�u�u�x�0�-����KĹ����^	�����0�&�u�x�w�}��������9��h�����%�:�u�u�%�>����	������D�����
��&�f�1�0�E���	����l��F1��*���
�&�
�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ǹ��^9��G�����u�u�u�u�w�}�WϹ�	����T��T��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�/�(���A�ѓ�VF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���T��Q��G݊�e�i�u�!��2����������^�����0�}��-��$����&����S��B�\��_�u�u�x�w�/�(���A�֓�VF��D��U���6�&�{�x�]�}�W���&���� V��R1�����
�'�6�o�'�2��������F��h��*���$��
�!��.�(������T9��R��!���a�3�8�f�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U���%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}����	����@��X	��*���u�%�&�2�4�8�(���
�ғ�@��G��U���;�_�u�u�w�}�W�������l^��h��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�:����&����P�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���Y�����h��M���%�u�h�&�3�1��������AN��D��]���;�1�<�
���8���HŹ��A��[�\��|�n�_�u�w���������\��h_��*���d�l�
�g�k�}��������E��X�����;�1�<�
�>���������A��^�U���;�<�;�1�6�����&����O�=N��U���9�
�:�
�8�-�C���
����V��h�I���!�%�3�
�d��Fϱ�Y����\��h��*���_�u�u��/�����&�Г�l ��\�*��i�u�!�
�8�4�(�������]��Y�����0�g�
� �f�j�(��Y�ƹ�@��R
�����9�b�3�
�e�d����B�����O=�����
�
� �d�b��E��Y����_	��T1�����}�;�<�;�3�3� ���O����
R��G]��Xʠ�&�2�0�}�2���������9��G�U���;�"�0�d��(�N���	���l�N��Uʥ�b��g�<��4�W����ο�_9��G1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N��*݊�
�a�<�
�>�f�W�������_W��Q��Mۊ�f�i�u�u�w�}�Wϰ�����l ��[�����=�;�}�'�4�3�(���A�ד�N��S��D���0�&�u�u�w�}�Wϰ�����l ��X����u�u�;�"�2�l�(���@�ߓ� F�d��U���u�;�"�0�n�;�(��&����[�������g�3�
�d��o�G���Y�����RNךU���u�u�0��;�m����Nƹ��l�N�����d�
� �l�`�-�W��s���F�Y����
� �l�d�'�}����Q����\��h��L���%�}�|�h�p�z�W������F�N�����d�
� �l�n�-�L���Yӈ��`��1��*��b�%�u�h�]�}�W���Y����a��~1�����<�u�=�;��8�(���Hʹ��lW��1��]���h�r�r�u�;�8�}���Y���C9��e��<��
�;�&�2�]�}�W���*����l ��_�*��i�u�u�u�w�}����+����lW��^ �����=�;�}�0��0�F؁�����
9��^��H��r�u�9�0�]�}�W���Y����a��~1�����<�n�u�u�9�*���&����U��G]��H�ߊu�u�u�u������&Ĺ��l�������0�
�8�d��(�F��&���F�_��U���0�_�u�u�w�}�(߁�����9��h��N���u�;�"�0�f����M����Z�=N��U���u�
�
�4���(���
����[����*���d�
� �d�a��E��Y���O��[�����u�u�u�
��<�6���L����@��=N��U����9�m�3��l�N���Y���F�N�����0�d�
� �f�m�(������	��T��M���
�d�f�%��t�J���^�Ʃ�@�N��U���;�"�0�d��(�F��&����F�Y����
� �d�c��n�K���Y���F��R�����3�
�d�d�'�}����Q����\��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����9�b�3�
�f�n���Y����V��[_�� ��b�%�u�h�]�}�W���Y����a��~1�*���&�2�"�0�w�.����	˹��l^��h�E���u�d�|�0�$�}�W���Y����lV��V��*Ҋ�;�&�2�_�w�}�����֓�F9�� _��F��u�u�u�u�w�3� ���H˹��lW��1��U���;�}�'�6�9�h����H�ѓ�N��S��D���0�&�u�u�w�}�Wϰ�����
9��h_�F���n�u�u�;� �8�Eށ�����
9��R�����u�u�u�
���(���
����[����*���d�
� �d�g��E��Y���O��[�����u�u�u�
���D���&����9F� ��&���g�3�
�d�b�-�W��s���F�G1��7��
�;�&�2� �8�Wǭ�����Q��B1�Mӊ�g�e�u�u�f�t����Y���F���*���
�;�&�2�]�}�W���*����l ��_�*��i�u�u�u�w�}����;�ѓ�]9��PN�����&�9�!�%�b�;�(��N����O�I�\ʰ�&�u�u�u�w�}����;�ӓ�]9��PUךU���0��9�a�1��F���	���l�N��Uʥ�b��f�<��4�W����ο�_9��G_�����e�`�%�}�~�`�P���Y����l�N��Uʥ�b��d�
�9�.��ԜY�Ƣ�D5��[�� ��e�
�f�i�w�}�W���Yӈ��`��1��*��l�%�u�=�9�u�����ޓ�F9��]��G��u�u�d�|�2�.�W���Y�����d��G���
�d�`�%�l�}�Wϰ�����9��h_�D���u�h�_�u�w�}�W���*����l ��_�*��"�0�u�:��2�ہ�����9��^��H��r�u�9�0�]�}�W���Y����V
��h��D��
�f�_�u�w�8�$���N����T��h�I���u�u�u�u�9�*���&����V��G]�����}�'�6�;�b�;�(��N����O�I�\ʰ�&�u�u�u�w�}��������U��_����u�u�;�"�2�o����Iʹ��Z�=N��U���u�
�
�4���(���
����[����*���a�3�
�`��o�G���Y�����RNךU���u�u�
�
�6��(ہ�����l�N�����f�3�
�g��n�K���Y���F��h^�����
�
�;�&�0�*����
����^��B1�F���}�|�h�r�p�}����s���F�G1��'����d�
�;�$�:�}���Y����V
��Q��G݊�f�i�u�u�w�}�Wϰ�����U��[��Fʢ�0�u�:�
�8�9����@¹��V�
N��R���9�0�_�u�w�}�W���*����U��Y��F�ߊu�u�0��;����H����[�N��U���;�"�0�g�1��Gց�Jӑ��]F��E1�����3�
�d�
�e�m�W���H����_��=N��U���u�0��9��(�N���	��ƹF��R��܊� �l�l�%�w�`�}���Y���]��R�����g�
�f�"�2�}��������U��[��G��u�u�d�|�2�.�W���Y�����d��*���l�d�%�n�w�}�����ѓ�F9�� 1��U��_�u�u�u�w��(���&����Z��_��]���
�8�f�3��j�(��I���W����ߊu�u�u�u���(�������T]ǻN�����9�
� �l�d�-�W��s���F�G1��7��
�;�&�2� �8�Wǭ�����9��hV�*��e�u�u�d�~�8����Y���F��hY��*Ҋ�;�&�2�_�w�}����ʹ��l_��h�I���u�u�u�u�'�j�5�������TF��R �����!�%�
� �o�h����P���A�R��U���u�u�u�%�`��C���&����9F� ��&���3�
�m�
�d�a�W���Y�����h<��4���
�;�&�2� �8�Wǭ����� 9��hV�*��e�u�u�d�~�8����Y���F��h^�����
�g�<�
�>�f�W�������]��Q��Eي�g�i�u�&�;�)�ׁ�����l��X�����8�c�3�
�a��E��Y����A9��Y
�����d�
�g�i�w�.����	ǹ��l^��h����0�
�8�g�1��Cց�K��ƹF��E1�����3�
�f�
�e�a�WǱ�&����l ��W�����'�:�
�:�3����J����l�N��*���1�
� �d�d��E��Yە��l��[�� ��b�
�g�:�w�8�(���Hǹ��lW��1��\�ߊu�u�'�6�9�h����H�ѓ�F�F��*���1�
� �d�f��Eϱ�Y����\��h��D��
�g�n�u�w�2�(���˹��lW��1��U��}�0�
�8�f����I¹��	��D�����m�3�
�e�b�-�^�ԜY�ƣ�l��SW�� ��g�
�g�i�w�.����	�ѓ�F9��W��Gʺ�u�0�
�8�f����A����]ǻN�����;�
� �m�f�-�W��Q����G��h��M���%�u�'�&�;�)�ށ�����l��dךU���x�%�e�� ��G���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l4��v'��*���#�1�<�
�>���������PF��G�����%�e��"��m��������lV��V��*ڊ�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��e��<���4�
�9�|�w�5��ԜY���F�N��E���"��e�4��1�(���
���F��1�����e�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
�6��(߁�	����l��D��I���
�
�4�����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4���(���
����@��YN�����&�u�x�u�w�-�G�������l��D�����2�
�'�6�m�-����
ۖ��l4��v'��Yʥ�e��"��g�-���	�֓�R��h^�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����+����lV��G1�����!�0�u�u�w�}�W���YӖ��l4��v'��*���&�2�i�u������&��ƹF�N�����_�u�u�u�w�}�W���&����z9��^ �����h�%�e�� ��G�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�4��
�g�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I����r/��1��*���
�;�&�2�6�.���������T��]���
�4��
�g�<�(���UӖ��l4��v'��E���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lV��V��*���4�
�9�|�w�5��ԜY���F�N��E���"��d�
�'�+����&����[��h^�����
�e�4�
�;�f�W���Y����_��=N��U���u�u�u�
��<�6���I����E
��^ �����h�%�e�� ��F߁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<�6���I����@��V�����'�6�&�{�z�W�W���&ù��D'��^�����2�4�&�2��/���	����@��h^�����
�e�u�
��<�6���I����TJ��h^�����
�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��e��<��
�%�#�1�~�)����Y���F�N��*ڊ�4��
�e�>�����DӖ��l4��v'��E�ߊu�u�u�u�;�8�}���Y���F�G1��'����d�
�;�$�:�K���&ù��D'��^�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(߁�����W��G1�����
�<�u�&�>�3�������KǻN��*ڊ�4��
�d�6���������l��^	�����u�u�'�6�$�u�(߁�����W��G1�����
�
�4���l��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�4���F���&����F��R ��U���u�u�u�u�'�m�%���0����R��[
�����2�i�u�
��<�6���H����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��@/��Dۊ�%�#�1�<��4�W��	�֓�R��h_�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��@/��Dۊ�;�&�2�4�$�:�W�������K��N������"��d��3��������]9��X��U���6�&�}�
��<�6���H�Ƽ�9��@/��Dۊ�'�2�u�
��<�6���H����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�e�� ��Fށ�	����O��_�����u�u�u�u�w��(���8����l��D��I���
�
�4���l�}���Y���V
��d��U���u�u�u�%�g�� ���H¹��l��R������"��d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��'����d�
�%�!�9�����ƭ�@�������{�x�_�u�w��(���8����l��A�����<�
�&�<�9�-����Y����V��G1��'����d�
�%�!�9�W���&����z9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��D'��\�����1�|�!�0�w�}�W���Y�����h<��4���g�4�
�9��3����E�Ƽ�9��@/��D؊�%�#�1�_�w�}�W������F�N��U���%�e��"��l�(�������]9��PN�U���
�4��
�e�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�e��"��l�(���
����@��YN�����&�u�x�u�w�-�G�������9��h��*���<�;�%�:�w�}����
�μ�9��@/��D���%�e��"��l�(����Ƽ�9��@/��D؊�%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�֓�R��h_�����9�|�u�=�9�W�W���Y���F��1�����d�
�;�&�0�a�W���&����z9��d��U���u�0�&�u�w�}�W���Y����lV��V��*���<�
�<�u�j�-�G�������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g�� ���H����l��h�����4�&�2�u�%�>���T���F��1�����d�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�g�� ���H����l��N��E���"��d�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N������"��d��-����PӒ��]FǻN��U���u�u�
�
�6��(�������W9��h��U��%�e��"��l�(�������F�N�����u�u�u�u�w�}�WϮ�I����r/��1��*���
�;�&�2�k�}�(߁�����U��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�I����r/��1��*���u�&�<�;�'�2����Y��ƹF��h^�����
�f�<�
�>���������PF��G�����%�e��"��l�[Ϯ�I����r/��1�����%�e��"��l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�4��
�d�<�(���P�Ƹ�V�N��U���u�u�%�e��*�>��&����Z�
N��E���"��d�n�w�}�W�������9F�N��U���u�
�
�4���D���&����[��h^�����
�f�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lV��V��*���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e��*�>��&����_��Y1�����&�2�
�'�4�g��������lV��V��*���4�
�9�y�'�m�%���0����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G�������9��h��\���=�;�_�u�w�}�W���Y����a��~1�*���#�1�<�
�>�}�JϮ�I����r/��1��*���n�u�u�u�w�8����Y���F�N��*ڊ�4��
�a�6���������Z�G1��'����d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�4��
�a�>�����
������T��[���_�u�u�
��<�6���M����@��V�����'�6�o�%�8�8�Ǯ�I����r/��B��*ڊ�4��
�a�'�8�[Ϯ�I����r/��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(߁�����R��G1�����!�0�u�u�w�}�W���YӖ��l4��v'��A���
�<�u�h�'�m�%���0����9F�N��U���0�_�u�u�w�}�W���&ù��D'��Z�����2�i�u�
��<�6���M����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�4���B���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l4��v'��@���
�9�
�;�$�:��������\������}�
�
�4���B���&������h<��4���`�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h^�����
�`�4�
�;�t�W������F�N��Uʥ�e��"��f���������@��S��*ڊ�4��
�`�6����Y���F��[�����u�u�u�u�w��(���8����l��A�����<�u�h�%�g�� ���Hƹ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���8����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��@/��Dߊ�;�&�2�4�$�:�(�������A	��D��*ڊ�4��
�`�w��(���8����l��PB��*ڊ�4��
�`�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��'����d�
�%�!�9�^Ϫ���ƹF�N��U���
�
�4���h���������h<��4���`�_�u�u�w�}����s���F�N������"��d��3����E�Ƽ�9��@/��Dߊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��D'��1��*���
�;�&�2�6�.��������@H�d��Uʥ�e��"��f�<�(���&����Z��D�����:�u�u�'�4�.�_���&����z9��V�����%�e��"��l��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�4���(��������YNךU���u�u�u�u������&¹��l��h�����i�u�
�
�6��(ށ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�֓�R��h_�����1�<�
�<�w�`����+����lW��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�I����r/��h�����4�&�2�u�%�>���T���F��1�����d�<�
�<��.����	����	F��X��¥�e��"��f�}�(߁�����9��R	�����"��d�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��'����d�4�
�;�t�W������F�N��Uʥ�e��"��f�4�(���Y����lV��V��*��u�u�u�u�2�.�W���Y���F���*����
�
�;�$�:�K���&ù��D'��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�G�������l��A�����<�u�&�<�9�-����
���9F���*����
�
�%�!�9��������@��h����%�:�0�&�'�m�%���0�ԓ�C9��SB��*ڊ�4��
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N������"��g�6�����Y����l�N��U���u�%�e�� ��E���&����Z��^	��Hʥ�e��"��e�<�(���B���F����ߊu�u�u�u�w�}�(߁�����9��h��*���&�2�i�u������&����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���8����Z��^	�����;�%�:�0�$�}�Z���YӖ��l4��v'��*���&�2�4�&�0�����CӖ��P����*����
�y�%�g�� ���K����TJ��h^�����
�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lV��V��*؊�%�#�1�|�#�8�W���Y���F���*����
�
�;�$�:�K���&ù��D'��UךU���u�u�9�0�]�}�W���Y���C9��e��<���<�
�<�u�j�-�G�������l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��<�6���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e��<���4�
�9�
�9�.����
����C��T�����&�}�
�
�6��(܁�	����F��1�����f�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h^�����
�
�%�#�3�t����Y���F�N��U���
�4��
��-��������TF���*����
�
�%�!�9�}���Y���V
��d��U���u�u�u�%�g�� ���J����E
��^ �����h�%�e�� ��D���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e��*�>�������TF��D��U���6�&�{�x�]�}�W���&����z9��^ �����&�<�;�%�8�}�W�������C9��e��<��u�
�
�4���(����Ƽ�9��@/��F���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��D'��1��*���|�u�=�;�]�}�W���Y���C9��e��<���<�
�<�u�j�-�G�������l�N��Uʰ�&�u�u�u�w�}�W���	�֓�R��h]�����2�i�u�
��<�6���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�e��"��i��������l�������%�:�0�&�w�p�W���	�֓�R��hZ�����1�<�
�<��.����	����	F��X��¥�e��"��c�<�(���UӖ��l4��v'��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��@/��A���
�9�|�u�?�3�}���Y���F�G1��'����a�4�
�;��������C9��e��<���4�
�9�n�w�}�W�������9F�N��U���u�
�
�4���(�������]9��PN�U���
�4��
��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�4�������Ӈ��Z��G�����u�x�u�u�'�m�%���0�ғ�]9��P1�����
�'�6�o�'�2����	�֓�R��hZ�����"��a�'�8�[Ϯ�I����r/��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G�������l��A��\ʡ�0�u�u�u�w�}�W���	�֓�R��hZ�����2�i�u�
��<�6���B���F����ߊu�u�u�u�w�}�(߁�����9��h��U��%�e��"��i����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�4��
�
�'�+����&����R��P �����&�{�x�_�w�}�(߁�����9��h��*���&�2�4�&�0�����CӖ��P����*����
�
�%�!�9�W���&����z9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�I����r/��h�����|�!�0�u�w�}�W���Y����lV��V��*ߊ�%�#�1�<��4�W��	�֓�R��h[�����1�_�u�u�w�}����s���F�N������"��`�6���������Z�G1��'����`�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��E���"��`�<��4�W�������A	��D�X�ߊu�u�
�
�6��(ځ�����l��^	�����u�u�'�6�$�u�(߁�����J��h^�����
�
�'�2�w��(���8����R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��<�6���&����_����ߊu�u�u�u�w�}�(߁�����9��h��U��%�e��"��h�}���Y���V
��d��U���u�u�u�%�g�� ���L����@��S��*ڊ�4��
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�����c�4�
�9��3��������]F��X�����x�u�u�%�g�� ���O����E
��^ �����&�<�;�%�8�}�W�������C9��e��<���4�
�9�y�'�m�%���0�Г�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���8����R��[
��U���;�_�u�u�w�}�W���&ù��D'��1��*���
�;�&�2�k�}�(߁�����9��h��N���u�u�u�0�$�}�W���Y���F��h^�����
�
�%�#�3�4�(���Y����lV��V��*܊�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h<��4���
�;�&�2�6�.��������@H�d��Uʥ�e��"��a�4�(���&����T��E��Oʥ�:�0�&�%�g�� ���O�Ƽ�9��@/��C���0�y�%�e��*�>�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e��"��k�������G��d��U���u�u�u�%�g�� ���O����@��S��*ڊ�4��
�n�w�}�W�������9F�N��U���u�
�
�4���(���
���F��1�����c�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l4��v'��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�4���(�������]9��P1�����
�'�6�o�'�2����	�֓�R��hY�����1�u�
�
�6��(؁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�e��*�>�������WO�C��U���u�u�u�u�w�-�G�������l��A�����<�u�h�%�g�� ���N����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��@/��B���
�9�
�;�$�:�K���&ù��D'�� 1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����a��~1�����<�u�&�<�9�-����
���9F���*����
�
�;�$�:��������\������}�
�
�4���[Ϯ�I����r/��h�����
�
�4����������F��P��U���u�u�<�u��-��������Z��S��*ڊ�4��
�
�'�+��������9F�N��U���u�
�
�4���(���
���F��1�����b�_�u�u�w�}����s���F�N������"��b�>�����DӖ��l4��v'��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����z9��V�����;�&�2�4�$�:�W�������K��N������"��m�6���������l��^	�����u�u�'�6�$�u�(߁�����9��h��Yʥ�e��"��o�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�4�����������[��=N��U���u�u�u�
��<�6���&����_��Y1����u�
�
�4���(�������F�N�����u�u�u�u�w�}�WϮ�I����r/��h�����<�
�<�u�j�-�G�������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����+����l^��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��e��<���<�
�<�
�$�4��������C��R������"��m�w��(���8����C��N��E���"��m�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����m�4�
�9�~�}����s���F�N������"��m�>�����DӖ��l4��v'��N���u�u�u�0�$�}�W���Y���F��h^�����
�
�;�&�0�a�W���&����z9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�%���0�ߓ�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h^�����
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�g�� ���@����E
����*����
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��E���"��l�4��1�^������F�N��U���%�e��"��d��������l��R������"��l�6����Y���F��[�����u�u�u�u�w��(���8����R��[
�����2�i�u�
��<�6���&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u������&ʹ��l�������%�:�0�&�w�p�W���	�֓�R��hW�����2�4�&�2��/���	����@��h^�����
�y�%�e��*�>���	������h<��4���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��v'��*���#�1�|�!�2�}�W���Y���F��h^�����
�
�;�&�0�a�W���&����z9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��@/��L���
�<�u�h�'�m�%���0�ߓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�6�9�3��G��Y����9��1��N�ߊu�u�x�%�c�����8����R��[
�����;�%�:�0�$�}�Z���YӖ��l5��[��<���4�
�9�
�$�4��������C��R�����0�u�%�&�0�>����-����l ��hX��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���=�;�_�u�w�}�W���Y����`��R
��*ڊ�%�#�1�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����lR��T�����e�4�
�9�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�
�
�4�1����H���R��1�G���n�u�u�%�c�����8����Z�V��E��g�$�n�_�w�}�ZϮ�M����_��~1�*���#�1�4�&�0�}����
���l�N��A���4�0��
�g�<�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�f�t�W������F�N��Uʥ�a��4�0���G���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�%�a��6�8�6���I����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�9��V��4���d�i�u�'���G݁�H��ƹF�N��A���4�0��
�f�<�(���Y����T��E�����x�_�u�u����������9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}�(ہ�����r/��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ǹ��R
��v'��D���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�6�9�3��F���DӇ��lV��\��E�ߠu�u�x�u����������9��h��U���<�;�%�:�2�.�W��Y����lR��T�����d�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�!�2�}�W���Y���F��hZ�����1��d�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*ފ�6�9�1��f��������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����*����W'��]��Hʴ�,�e�c�g�&�f�}���Y����lR��T�����d�
�%�#�3�<����Y����V��C�U���%�a��4�2��(�������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�f�3�:�l�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��P�Ƹ�V�N��U���u�u�%�a��<����&�Փ�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�i�$�������U��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1��&���0��
�a�k�}����&����BV��=N��U���%�a��4�2��(�������WF��D��U���6�&�{�x�]�}�W���&����V��h_�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���Hǹ��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�_�u�w�}�W���Y����`��R
��*���4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��d�����
�a�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
��>����0����[��E��*��
�d�_�u�w�p�W���&����V��h_�����9�u�&�<�9�-����
���9F���*���9�1��d��-��������]9��X��U���6�&�}�%�4�q��������V��c1��Dފ�&�
�f�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���a�3�8�d�~�t����Y���F�N��U���
�6�9�1��l�(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�6�;�9�>��&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h=������d�4�
�;�}����Ӗ��P��N����u�
�
�6�;�9�>�������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�b�3�:�k�^������F�N��U���%�a��4�2��(ށ�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�4�1����H����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�9��V��4���u�h�4�,�g�k�E���B���F���*���9�1��g�6�����
������T��[���_�u�u�
��>����0�ԓ�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!��.�(���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�o�;���P�Ƹ�V�N��U���u�u�%�a��<����&����l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u����������l��A��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��1������
�u�h�6�$�G��K����9l�N�U���
�6�9�1��n�����ƭ�@�������{�x�_�u�w��(�������lU��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�(���&��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�O������F��R ��U���u�u�u�u�'�i�$������� 9��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}�(ہ�����r/��h�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N��A���4�0��
�w�`����I����l��=d��U���u�
�
�6�;�9�>�������WF��D��U���6�&�{�x�]�}�W���&����V��hZ�����1�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���&����OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���@����l^�N�����u�u�u�u�w�}����*����W'��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ǹ��R
��v'��*���#�1�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʥ�a��4�0���W������lP��h����u�x�u�
��>����0�ӓ�C9��SN�����u�'�6�&�y�p�}���Y����`��R
��*ߊ�%�#�1�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��hV��\ʡ�0�u�u�u�w�}�W���	�ғ�P��S/��@���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��V��4���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�a��6�8�6���Y����A��hX�*��_�u�u�x�w��(�������lP��G1��ʴ�&�2�u�'�4�.�Y��s���C9��d�����
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��^�����|�|�!�0�w�}�W���Y�����h=������c�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1��&���0��
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�i�$�������F���*ڊ�e�
�d�_�w�}�Z���&ǹ��R
��v'��*���#�1�4�&�0�}����
���l�N��A���4�0��
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��Dڊ�&�
�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�~�)����Y���F�N��*ފ�6�9�1��`�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�a��4�0���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�M����_��~1�I���'�
�
�e��m�}���Y���C9��d�����
�
�%�#�3�<����Y����V��C�U���%�a��4�2��(ׁ�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�d�
�&��m�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�d�1�0�F���PӒ��]FǻN��U���u�u�
�
�4�1����A����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�c�����8����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h=������l�i�u�%��(��&����9F�C�����4�0�������Ӈ��Z��G�����u�x�u�u�'�i�$�������
9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O����ߊu�u�u�u�w�}�(ہ�����r/��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�M����_��~1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hY��*ڊ�%�#�1�u���(߁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�b��m�������G��d��U���u�u�u�%�`��G���&����Z��^	��Hʥ�b��e�4��1�L���Y�����RNךU���u�u�u�u���(߁�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�b��g�4�(���&����T��E��Oʥ�:�0�&�%�`��G���&Ĺ��9��R	�����e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��u1�����9�|�u�=�9�W�W���Y���F�� 1��E���
�<�u�h�'�j�5��s���F�R��U���u�u�u�u�w�-�@���I����@��S��*݊�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��^�����1�<�
�<�w�.����	����@�CךU���
�
�
�e�6���������l��^	�����u�u�'�6�$�u�(؁�&�֓�C9��SB��*݊�
�e�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���e�4�
�9�~�}����s���F�N������d�
�%�!�9���������h,��E���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�e�6���������Z�G1��7��
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�e�<��4�(�������A	��N�����&�%�b��f�q����;����C��N��B���d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lQ��h_�����9�|�u�=�9�W�W���Y���F�� 1��Dڊ�;�&�2�i�w��(���I���F�N�����u�u�u�u�w�}����;����Z��^	��Hʥ�b��d�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F�� 1��Dۊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��l��������l��h�����%�:�u�u�%�>����&Ĺ��W��G1�����
�
�
�d�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�d�4��1�^������F�N��U���%�b��d��-��������TF���*���d�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
��l��������l��R������d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�d�<�
�>�}����Ӗ��P��N����u�
�
�
�f�4�(���&����T��E��Oʥ�:�0�&�%�`��F��	�ѓ�lW��G��Yʥ�b��d�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*���4�
�9�|�w�5��ԜY���F�N��B���d�
�;�&�0�a�W���&����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lW��^ �����h�%�b��f�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���d�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(�������W9��h��*���<�;�%�:�w�}����
�μ�9��\�����1�u�
�
��o��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�e�<�(���P�Ƹ�V�N��U���u�u�%�b��l�(�������]9��PN�U���
�
�g�4��1�L���Y�����RNךU���u�u�u�u���(�������W9��h��U��%�b��d��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�
�g�>�����
������T��[���_�u�u�
���E���&����R��P �����o�%�:�0�$�-�@���H����lQ��h_�����y�%�b��f��������F��P��U���u�u�<�u��-��������Z��S��*݊�
�g�4�
�;�t�W������F�N��Uʥ�b��d�
�9�.���Y����q9��d��U���u�0�&�u�w�}�W���Y����lQ��h_�����<�u�h�%�`��F݁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b��d�
�'�+����&����R��P �����&�{�x�_�w�}�(؁�&�Փ�C9��S1��*���
�&�<�;�'�2�W�������@N�� 1��Dي�%�#�1�u���(�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
���D���&����F��R ��U���u�u�u�u�'�j�5��&����_��Y1����u�
�
�
�d�<�(���B���F����ߊu�u�u�u�w�}�(؁�&�Փ�C9��S1��*���u�h�%�b��l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
��n�����ƭ�@�������{�x�_�u�w��(���J����@��V�����'�6�o�%�8�8�Ǯ�N���� J��hY��*���%�0�y�%�`��F܁�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�f�6�����Y����l�N��U���u�%�b��f��������C9��u1�N���u�u�u�0�$�}�W���Y���F��hY��*���<�
�<�u�j�-�@���H����V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�b��f���������@��V�����'�6�&�{�z�W�W���&Ĺ��R��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B���d�
�%�#�3�}�(؁�&�ғ�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���M����E
��N�����u�u�u�u�w�}����;����R��[
�����2�i�u�
���C���&����9F�N��U���0�_�u�u�w�}�W���&Ĺ��R��G1�����
�<�u�h�'�j�5��&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(�������TF��D��U���6�&�{�x�]�}�W���&����l��D�����2�
�'�6�m�-����
ۖ��l$��B��*݊�
�a�%�0�{�-�@���Hǹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��i�������G��d��U���u�u�u�%�`��Fہ�����Z�G1��7��n�u�u�u�w�8����Y���F�N��*݊�
�a�<�
�>�}�JϮ�N����9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`��Fځ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��[�����1�<�
�<��.����	����	F��X��¥�b��d�
�'�+����&Ĺ��S��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����l��A��\ʡ�0�u�u�u�w�}�W���	�ѓ�lW��V�����;�&�2�i�w��(���L����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��[�����1�<�
�<�w�`����;����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(؁�&�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����q9��h�����4�&�2�
�%�>�MϮ�������h,��@���
�
�
�`�'�8�[Ϯ�N����9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(�������WO�C��U���u�u�u�u�w�-�@���Hƹ��l��R������d�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�`�>�����DӖ��l$��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@���H����E
��^ �����&�<�;�%�8�8����T�����h,��*���#�1�<�
�>���������PF��G�����%�b��d�6����	�ѓ�lW��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&Ĺ��9��h��*���&�2�i�u���(ށ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lW��G1�����
�<�u�h�'�j�5�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`��F���&����R��P �����&�{�x�_�w�}�(؁�&¹��l��h�����%�:�u�u�%�>����&Ĺ��J��hY��*ۊ�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����q9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���u�h�%�b��l����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(݁�	����l��D�����2�
�'�6�m�-����
ۖ��l$��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b��g�4��1�^������F�N��U���%�b��g�6���������Z�G1��7���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*؊�;�&�2�4�$�:�W�������K��N������g�<�
�>���������PF��G�����%�b��g�w��(���&����F�� 1��G���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��9��h��\���=�;�_�u�w�}�W���Y����q9��^ �����h�%�b��e�W�W���Y�Ʃ�@�N��U���u�u�%�b��o���������h,��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1��7���4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ѓ�lU��G1�����!�0�u�u�w�}�W���YӖ��l$��h�����<�
�<�u�j�-�@���J����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���
�;�&�2�k�}�(؁�&����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�N����l��D�����2�
�'�6�m�-����
ۖ��l$��N��B���f�%�0�y�'�j�5�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��f�6�����Y����l�N��U���u�%�b��d�4�(���Y����lQ��h]�U���u�u�0�&�w�}�W���Y�����h,��*���&�2�i�u���(܁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b��a�4��1�(���
����@��YN�����&�u�x�u�w�-�@���M����E
��^ �����&�<�;�%�8�}�W�������C9��u1�����9�y�%�b��i��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*݊�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�b��i��������l��R������a�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���a�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q����;�ғ�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l$��h�����|�!�0�u�w�}�W���Y����lQ��hZ�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ہ�����Z�G1��7���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�lS��G1�����
�<�u�&�>�3�������KǻN��*݊�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�`��B���&������h,��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��1��*���|�u�=�;�]�}�W���Y���C9��u1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h,��*���#�1�<�
�>�}�JϮ�N����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����;�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����q9��^ �����&�<�;�%�8�}�W�������C9��u1�U���
�
�
�'�0�}�(؁�&ƹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F�� 1��@�ߊu�u�u�u�;�8�}���Y���F�G1��7���<�
�<�u�j�-�@���L����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hY��*܊�%�#�1�u���(ف�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�b��k�������G��d��U���u�u�u�%�`��A���&����Z��^	��Hʥ�b��c�4��1�L���Y�����RNךU���u�u�u�u���(ف�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�b��a�4�(���&����T��E��Oʥ�:�0�&�%�`��A���&Ĺ��9��R	�����c�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��u1�����9�|�u�=�9�W�W���Y���F�� 1��C���
�<�u�h�'�j�5��s���F�R��U���u�u�u�u�w�-�@���O����@��S��*݊�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9�� 1��*���
�;�&�2�6�.��������@H�d��Uʥ�b��b�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1��7���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h,��*���#�1�|�!�2�}�W���Y���F��hY��*݊�%�#�1�<��4�W��	�ѓ�lQ��G1���ߊu�u�u�u�;�8�}���Y���F�G1��7���4�
�9�
�9�.���Y����q9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&Ĺ��9��h��U���<�;�%�:�2�.�W��Y����lQ��hY�����2�4�&�2��/���	����@��hY��*���%�b��b�'�8�[Ϯ�N����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`��@���&����F��R ��U���u�u�u�u�'�j�5�������TF���*���n�u�u�u�w�8����Y���F�N��*݊�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b��e��������l�������%�:�0�&�w�p�W���	�ѓ�l^��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B���m�4�
�9�{�-�@���A����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(ׁ�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�@���A����E
��^ �����h�%�b��o�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b��m�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l$��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*Ҋ�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(؁�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�b��m�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h,��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.����;�ߓ�C9��SB��*݊�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��7���4�
�9�|�w�5��ԜY���F�N��B���l�4�
�9��3����E�Ƽ�9��1��*���n�u�u�u�w�8����Y���F�N��*݊�
�
�%�#�3�4�(���Y����lQ��hW�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l$��h�����4�&�2�u�%�>���T���F�� 1��L���
�<�
�&�>�3����Y�Ƽ�\��DF��B���l�u�
�
������Y����q9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(؁�&ʹ��l��R������l�_�u�w�}�W������F�N��Uʥ�b��l�<��4�W��	�ѓ�l_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(߁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�N���I����E
��N�����u�u�u�u�w�}����4�֓�C9��S1��*���u�h�%�l��m������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�d�:�������T9��D��*���6�o�%�:�2�.����4���C9��z1�����y�%�l��g�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��L���e�4�
�9�~�}����s���F�N������e�<�
�>�}�JϮ�@����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�lV��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��8��
�%�#�1�>�����
������T��[���_�u�u�
���G���&����Z��^	�����;�%�:�u�w�/����Q����~9��h�����u�
�
�
�g�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�e�6�����Y����l�N��U���u�%�l��f���������@��S��*ӊ�
�e�4�
�;�f�W���Y����_��=N��U���u�u�u�
���G���&����Z��^	��Hʥ�l��d�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�e�<��4�W�������A	��D�X�ߊu�u�
�
��m��������@��h����%�:�0�&�'�d�:��UӖ��l+��1�����%�l��d��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���e�4�
�9�~�}����s���F�N������d�
�;�$�:�K���&ʹ��V��N��U���0�&�u�u�w�}�W���YӖ��l+��1��*���u�h�%�l��l�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����d�
�%�!�9�����ƭ�@�������{�x�_�u�w��(���H����E
��^ �����&�<�;�%�8�}�W�������C9��z1�*���#�1�u�
���F���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��l�������G��d��U���u�u�u�%�n��Fށ�	����l��D��I���
�
�
�d�6����Y���F��[�����u�u�u�u�w��(���H����E
��^ �����h�%�l��f���������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
�f�4�(���Y����T��E�����x�_�u�u���(�������T9��D��*���6�o�%�:�2�.����4������h#��D���0�y�%�l��l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�d�4��1�^������F�N��U���%�l��d��3����E�Ƽ�
9��_�U���u�u�0�&�w�}�W���Y�����h#��D���
�<�u�h�'�d�:��&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�l��d��-��������TF��D��U���6�&�{�x�]�}�W���&����l��A�����<�
�&�<�9�-����Y����V��G1��8��
�%�#�1�w��(���K����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(�������WO�C��U���u�u�u�u�w�-�N���H����l��h�����i�u�
�
��o������ƹF�N�����_�u�u�u�w�}�W���&����l��A�����<�u�h�%�n��F݁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
���E���&����R��P �����&�{�x�_�w�}�(ց�&�ԓ�]9��P1�����
�'�6�o�'�2����	�ߓ�lW����*���g�%�0�y�'�d�:��&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�e�<�(���P�Ƹ�V�N��U���u�u�%�l��l�(���
���F��1��D��u�u�u�u�2�.�W���Y���F���*���g�<�
�<�w�`����4����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�l��l�(�������]9��PN�����u�'�6�&�y�p�}���Y����~9��h�����<�
�<�
�$�4��������C��R������d�
�%�!�9�W���&����l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ց�&�Փ�C9��SG�����u�u�u�u�w�}�WϮ�@���� 9��h��*���&�2�i�u���(�������W]ǻN��U���9�0�_�u�w�}�W���Y����~9��h�����<�
�<�u�j�-�N���H����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���J����@��V�����'�6�&�{�z�W�W���&ʹ��U��Y1�����&�2�
�'�4�g��������l_��h_�U���
�
�f�%�2�q����4����R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
���D���&����F��R ��U���u�u�u�u�'�d�:��&����Z�
N��L���d�n�u�u�w�}����Y���F�N��U���
�
�f�<��4�W��	�ߓ�lW��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�:��&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��z1�*���#�1�<�
�>���������PF��G�����%�l��d��-����Y����~9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ʹ��R��G1�����!�0�u�u�w�}�W���YӖ��l+��1��*���
�;�&�2�k�}�(ց�&�ғ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��z1�*���#�1�<�
�>�}�JϮ�@����9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��Z�����2�4�&�2��/���	����@��hW��*��u�
�
�
�c�-���	�ߓ�lW��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���M����E
��N�����u�u�u�u�w�}����4����Z��^	��Hʥ�l��d�n�w�}�W�������9F�N��U���u�
�
�
�c�4�(���Y����l_��h_�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����4����R��[
�����2�4�&�2�w�/����W���F�G1��8��
�%�#�1�>�����
����l��TN����0�&�%�l��l�(������C9��z1�*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�
9��[�����1�|�!�0�w�}�W���Y�����h#��@���
�9�
�;�$�:�K���&ʹ��S��G1���ߊu�u�u�u�;�8�}���Y���F�G1��8��
�%�#�1�>�����DӖ��l+��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����~9��h�����4�&�2�u�%�>���T���F��1��Dߊ�;�&�2�4�$�:�(�������A	��D��*ӊ�
�`�u�
���B�������l_��h_�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����l��A��\ʡ�0�u�u�u�w�}�W���	�ߓ�lW��^ �����h�%�l��f�f�W���Y����_��=N��U���u�u�u�
���B���&����[��hW��*���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�lW��G1�����
�<�u�&�>�3�������KǻN��*ӊ�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�n��F���&������h#��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�
9��1��*���|�u�=�;�]�}�W���Y���C9��z1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h#��*���#�1�<�
�>�}�JϮ�@����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����4�ד�]9��PN�����u�'�6�&�y�p�}���Y����~9��^ �����&�<�;�%�8�}�W�������C9��z1�U���
�
�
�'�0�}�(ց�&¹��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F��1��D�ߊu�u�u�u�;�8�}���Y���F�G1��8���<�
�<�u�j�-�N���H����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hW��*؊�%�#�1�u���(݁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l��o�������G��d��U���u�u�u�%�n��E���&����Z��^	��Hʥ�l��g�4��1�L���Y�����RNךU���u�u�u�u���(݁�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�l��e�4�(���&����T��E��Oʥ�:�0�&�%�n��E���&ʹ��9��R	�����g�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��z1�����9�|�u�=�9�W�W���Y���F��1��G���
�<�u�h�'�d�:��s���F�R��U���u�u�u�u�w�-�N���K����@��S��*ӊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�l��f�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1��8���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h#��*���#�1�|�!�2�}�W���Y���F��hW��*ي�%�#�1�<��4�W��	�ߓ�lU��G1���ߊu�u�u�u�;�8�}���Y���F�G1��8���4�
�9�
�9�.���Y����~9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ʹ�� 9��h��U���<�;�%�:�2�.�W��Y����l_��h]�����2�4�&�2��/���	����@��hW��*���%�l��f�'�8�[Ϯ�@����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�n��D���&����F��R ��U���u�u�u�u�'�d�:�������TF���*���n�u�u�u�w�8����Y���F�N��*ӊ�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�l��i��������l�������%�:�0�&�w�p�W���	�ߓ�lR��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��L���a�4�
�9�{�-�N���M����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(ہ�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�N���M����E
��^ �����h�%�l��c�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�l��a�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l+��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hW��*ފ�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(ց�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�l��a�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h#��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.����4�ӓ�C9��SB��*ӊ�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��8���4�
�9�|�w�5��ԜY���F�N��L���`�4�
�9��3����E�Ƽ�
9��1��*���n�u�u�u�w�8����Y���F�N��*ӊ�
�
�%�#�3�4�(���Y����l_��h[�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l+��h�����4�&�2�u�%�>���T���F��1��@���
�<�
�&�>�3����Y�Ƽ�\��DF��L���`�u�
�
������Y����~9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(ց�&ƹ��l��R������`�_�u�w�}�W������F�N��Uʥ�l��`�<��4�W��	�ߓ�lS��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(ف�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�N���O����E
��N�����u�u�u�u�w�}����4�Г�C9��S1��*���u�h�%�l��k������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�d�:�������T9��D��*���6�o�%�:�2�.����4���C9��z1�����y�%�l��a�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��L���c�4�
�9�~�}����s���F�N������c�<�
�>�}�JϮ�@����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�lP��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��8���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�l��j��������l��h�����%�:�u�u�%�>����&ʹ��9��h��Yʥ�l��b�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ӊ�
�
�%�#�3�t����Y���F�N��U���
�
�
�%�!�9���������h#��*���#�1�_�u�w�}�W������F�N��Uʥ�l��b�4��1�(���
���F��1��B���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��z1�����<�u�&�<�9�-����
���9F���*���
�;�&�2�6�.���������T��]���
�
�y�%�n��@�������l_��hY�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����4�ѓ�C9��SG�����u�u�u�u�w�}�WϮ�@����l��D��I���
�
�
�n�w�}�W�������9F�N��U���u�
�
�
��3����E�Ƽ�
9�� 1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�N���A����E
��^ �����&�<�;�%�8�8����T�����h#��*���#�1�<�
�>���������PF��G�����%�l��m�6����	�ߓ�l^��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&ʹ��9��h��*���&�2�i�u���(ׁ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�l^��G1�����
�<�u�h�'�d�:�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n��O���&����R��P �����&�{�x�_�w�}�(ց�&˹��l��h�����%�:�u�u�%�>����&ʹ��J��hW��*Ҋ�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����~9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�
9��1��*���u�h�%�l��e����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ӊ�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(ց�	����l��D�����2�
�'�6�m�-����
ۖ��l+��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�l��l�4��1�^������F�N��U���%�l��l�6���������Z�G1��8���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hW��*ӊ�;�&�2�4�$�:�W�������K��N������l�<�
�>���������PF��G�����%�l��l�w��(���&����F��1��L���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ʹ��
9��h��\���=�;�_�u�w�}�W���Y����~9��^ �����h�%�l��n�W�W���Y�Ʃ�@�N��U���u�u�%�l��d���������h#��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�8�(���Hù��lW��1��U��_�u�u�u�w��(���&����Z��_��]���
�8�c�3��k�(��I���W����ߊu�u�u�u�2���������^��UךU���0�
�8�d��(�F��&���FǻN��U���
�
�
�e�>��������@��C��*���m�b�%�}�~�`�P���Y����l�N��Uʦ�9�!�%�e�1��G���	��ƹF��R����
� �d�f��n�K���Y���F��hW��*���<�
�<�u�?�3�_���&����l ��Y�����|�h�r�r�w�1��ԜY���F��[1�����3�
�e�g�'�f�W���
����^��h��D��
�g�i�u�f�}����Q����Z9��E1�����
�
�
� �f�h�(��DӇ��P	��C1��A��u�9�0�w�u�W�W�������CW��Q��E���%�u�h�w�u�*��������l ��h"�����d�&�3�
�g�d����Y����\��h��*���0�&�u�e�l�}�Wϭ�����S��B1�B݊�g�i�u�d�w�5����5����u	��{��*ފ�
�
� �d�b��E������]��[��B���9�0�w�w�]�}�W���&����9��h_�F���u�h�w�w� �8�WǷ�&����\��X��A���&�3�
�e�n�-�W���	����@��AZ��\ʰ�&�u�e�n�w�}��������l ��^�*��i�u�d�u�?�3�_�������A9��X��*ۊ�
� �d�`��o�JϿ�&����G9��1��U���0�w�w�_�w�}��������U��W�����h�w�w�"�2�}��������l*��G1��D���3�
�e�l�'�}�W�������l
��h*�����u�e�n�u�w�.����	�ߓ�F9��_��G��u�d�u�=�9�u�;���&����	��hZ��*��� �d�`�
�e�`��������_��G�����w�w�_�u�w�8�(���H����Q��G\��H���w�"�0�u�#�-����Jʹ��[��G1�����9�a��u�;�8�U���s���@��C��E���
�g�b�%�w�`�}���Y���C9��z1�����<�u�=�;��8�(���H����lW��1��]���h�r�r�u�;�8�}���Y���C9��z1�*���&�2�_�u�w�8�(���K¹��lW��1��U��_�u�u�u�w��(���&����Z��_��]���
�8�d�
�"�l�@ށ�K���F�G�����_�u�u�u�w�8�(���Kù��lW�� 1��N���u�&�9�!�'�o����K�֓� F�d��U���u�%�l��`�4�(���Y����N��[1�����3�
�e�b�'�u�^��^���V
��d��U���u�&�9�!�'�l����K�Փ� ]ǻN�����8�g�
� �f�i�(��E��ƹF�N��*ӊ�
�
�;�&�0�*����
����^��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�g�
� �f�i�(��s���@��C��A���
�g�a�%�w�`�}���Y���C9��z1�*���&�2�"�0�w�.����	�ѓ�F9��W��G��u�u�d�|�2�.�W���Y�����h��Gي� �d�a�
�d�W�W�������CT��Q��G���%�u�h�_�w�}�W���&ʹ��U��Y1��ʢ�0�u�&�9�#�-�O���&����l��G��U��|�0�&�u�w�}�W���
����^��h��D���
�f�_�u�w�8�(���K����R��G\��H���w�"�0�u�#�-����Jʹ��[��G1�����9�a�a�u�;�8�U���s���@��C��*���m�l�%�u�j��Uϩ�����^��B1�L���u�u�%�6�9�)����I�Ʃ�@�L�U���&�9�!�%��(�O���	���D�������8�
� �m�n�-�W���	����@��AZ��\ʰ�&�u�e�n�w�}��������U��^�����h�_�u�u�w�}�(ց�&����l�������0�
�8�
�"�e�D���Q���A��N�����u�u�u�u�'�d�:��&����Z��N�����!�%�
� �o�l����D������YN����� �m�l�%�w�}��������ER��N�����e�n�u�u�$�1����&����W��G]��H�ߊu�u�u�u���(ہ�������YN�����8�g�3�
�c��E��Y���O��[�����u�u�u�0��0�B���&����l��=N��U���
�8�m�3��k�(��E���F��R �����3�
�f�
�f�`��������_��vG�����w�w�_�u�w�8�(���@����V��h�I���u�u�u�u�'�d�:�������TF��R �����!�%�
� �o�h����P���A�R��U���u�u�u�&�;�)�؁�����9��d��Uʦ�9�!�%�3��i�(��E���F��R �����3�
�f�
�f�`��������_��G�����w�w�_�u�w�0�(ށ�����
9��R�����9�2�6�#�4�2�_�������]��Y�����<��'��8��(���&����P��UךU���8�
�
�
�"�l�G߁�H���@��[�����6�:�}�0�>�8��������Z*��^1�����:�
�
�
��8�(��N����O��N�����3�
�f�
�f�a�W�������A9��X��*���
�e�}�u�w�}�������9������