-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�g�d����}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e� �&�4�2��(���Y����g"��x)��*�����}�`�3�*����P���F��h��Oʜ�u��
���f�W���	�֓�]��[��<���4�
�9�u�w��$���5����l�N��E���&�4�0���}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��D�����
�
�%�#�3�g�>���-����t/��=N��U���
�;�6�9�3��E��0�Ɵ�w9��p'��#����u�d�u�8�3���B�����h;�����1��g�4��1�W���7ӵ��l*��~-�U���%�e� �&�6�8�6���Y�ƅ�5��h"��<������}�b�9� ���Y����F�G1�� ���4�0��
��-����Cӯ��`2��{!��6�ߊu�u�
�
�9�>����0���/��d:��9�������w�l�W������]ǻN��*ڊ�;�6�9�1��i��������z(��c*��:���n�u�u�%�g���������F��~ ��!�����
����_������\F��d��Uʥ�e� �&�4�2��(ځ�	����\��yN��1�����_�u�w��(�������r/��T��;ʆ�������8���H�ƨ�D��^����u�
�
�;�4�1����O����E
��N��U���
���n�w�}����,����_��~1�Oʜ�u��
����2���+������Y��E��u�u�%�e��.����8����R��[
��U��������W�W���&ù��@��R
��*���u������4���:����W��S�����|�_�u�u����������l^��G1�����u��
���L���YӖ��l3��T�����l�o��u���8���&����|4�[�����:�e�n�u�w�-�G���
����W'��1��*���u�u�����0���s���C9��b ������
�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I����P��S/��Dڊ�%�#�1�o��}�#���6����9F���*���6�9�1��f�}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��D�����
�d�4�
�;�}�W���*����|!��d��Uʥ�e� �&�4�2��(��Cӯ��`2��{!��6�����u�d�w�2����I��ƹF��h^�����9�1��d��-����Cӯ��`2��{!��6�ߊu�u�
�
�9�>����0����	F��=��*����
����u�BϺ�����O��N����� �&�4�0���D���&����	F��=��*����n�u�u�'�m�"�������z9��T��;ʆ�������8���H�ƨ�D��^����u�
�
�;�4�1����Hǹ��l��T��;ʆ�����]�}�W���&����R
��v'��@���u��
���(���-���S��X����n�u�u�%�g���������S��G1�����u��
���L���YӖ��l5��[��<��o������0���/����aF�N�����u�|�_�u�w��(�������lV��G1����������4�ԜY�Ƽ�9��V��4���u�u� �u���8���&����|4�_�����:�e�n�u�w�-�C�������z9��V�����u� �u����>��Y����lR��T�����g�o�����;���:����g)��]����!�u�|�_�w�}�(ہ�����r/��h�����o������0���s���C9��d�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}����*����W'��1��*���u�u� �u���8���B�����h=������a�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����V��hZ�����1�o�����;���:���F��1������
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�M����_��~1�����9�u�u� �w�	�(���0��ƹF��hZ�����1��c�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ǹ��R
��v'��*���#�1�o����3���>����F�G1��&���0��
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ғ�P��S/��B���
�9�u�u��}�#���6����9F���*���9�1��m�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����`��R
��*Ҋ�%�#�1�o��	�$���5����l�N��A���4�0��
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l5��[��<���4�
�9�u�w��W���&����p]ǻN��*ފ�6�9�1��f�}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lR��T�����d�
�%�#�3�g�8���*����|!��d��Uʥ�a��4�0���F��6����g"��x)��*�����}�d�3�*����P���F��1������
�d�4��1�W���,�Ɵ�w9��p'�����u�
�
�6�;�9�>��Y�ƃ�gF��s1��2������u�d�}�������9F���*���9�1��d��-����Cө��5��h"��<��u�u�%�a��<����&���)��=��*����
����u�FϺ�����O��N������4�0���n��������|3��d:��9����_�u�u����������F��x;��&���������W��Y����G	�UךU���
�
�6�9�3��Fہ�	����\��b:��!�����n�u�w�-�C�������z9��T�� ����
�����#���Q����\��XN�N���u�%�a��6�8�6���L����E
��N��!ʆ�����]�}�W���&����	F��=��*����
����u�BϺ�����O��N������e�4�
�;�}�W���*����|!��d��Uʥ�b��d�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�N����l��A��Oʜ�u��
���f�W���	�ѓ�lT�'��&���������W��Y����G	�UךU���
�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�
�w�}�9ύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����q9��V�����u������4�ԜY�Ƽ�9��N�<����
�����#���Q����\��XN�N���u�%�b��c�<�(���Y�ƅ�5��h"��<��u�u�%�b��h�Mϗ�Y����)��t1��6���u�d�u�:�9�2�G��Y����lQ��h[�����1�o��u���8���B�����h,��U���������!���6���F��@ ��U���_�u�u�
���(������/��d:��9����_�u�u���(���Y����g"��x)��*�����}�`�3�*����P���F�� 1��B���
�9�u�u���3���>����F�G1��7��o��u����>���<����N��
�����e�n�u�u�'�j�5�������WF��~ ��!�����n�u�w�-�@���@����}F��s1��2������u�f�}�������9F���*���
�%�#�1�m��W���&����p]ǻN��*݊�
�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����;����R��[
��U��������W�W���&Ĺ��W�'��&���������W��Y����G	�UךU���
�
�
�d�6�����Y����g"��x)��N���u�%�b��f�}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��\�����1�o��u���8���B�����h,��F���u��
���(���-���S��X����n�u�u�%�`��F܁�	����\��yN��1�����_�u�w��(���M����}F��s1��2������u�f�}�������9F���*���a�4�
�9�w�}�9ύ�=����z%��N������d�u�u���3���>����v%��eN��@ʱ�"�!�u�|�]�}�W���&����l��A��Oʜ�u��
���f�W���	�ߓ�lV�'��&���������W��Y����G	�UךU���
�
�
�
�'�+���0�Ɵ�w9��p'�����u�
�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����~9��V�����u������4�ԜY�Ƽ�
9��N�<����
�����#���Q����\��XN�N���u�%�l��e�<�(���Y�ƅ�5��h"��<��u�u�%�l��n�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����l_��h]�����1�o��u���8���B�����h#��U���������!���6���F��@ ��U���_�u�u�
���(������/��d:��9����_�u�u���(���Y����g"��x)��*�����}�d�3�*����P���F��1��@���
�9�u�u���3���>����F�G1��8��o��u����>���<����N��
�����e�n�u�u�'�d�:�������WF��~ ��!�����n�u�w�-�N���N����}F��s1��2������u�d�}�������9F���*���
�%�#�1�m��W���&����p]ǻN��*ӊ�
�u�u����;���:����g)��]����!�u�|�_�w�}�(ց�&˹��l��T��;ʆ�����]�}�W���&����	F��=��*����
����u�FϺ�����O��N������l�4�
�;�}�W���*����|!��d��Uʥ�l��d�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���&ʹ��V��G1�����u��
���L���YӖ��l+��N�<����
�����#���Q����\��XN�N���u�%�l��f���������}F��s1��2���_�u�u�
���E��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����h#��G���
�9�u�u���3���>����F�G1��8��u�u�����0���/����aF�N�����u�|�_�u�w��(���J����E
��N��U���
���n�w�}����4����	F��=��*����
����u�FϺ�����O��N������d�
�%�!�9�Mϗ�Y����)��tUךU���
�
�
�`�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ߓ�lW��V�����u������4���s����9l��E����� �0�7�=�!�2�W���K�Ԉ�r �������u�!�'�7�#�}�8���>����r2��y1��3���u����]�}�W�������VF��e+��0��������}�ϼ������_�����0�<�_�u�w�0�E��=ǧ��J��D1��*��a�a�.����"��� ����K��{=��;���
���h�{��(���,����k#��B��&�������j�>�������K��"��<�������e�s�G��I߮��l/��b:��'���:�=�'�y���.���5����V�V�EƝ������n�[���&����g6��Y��Y���
��
��j�q�;��� ����c[��"��&����h�a�`���$���5��� U��UךU���:�&�4�!�6�����&����P9��N��1�����o�u�f�f�W�������R��V�����
�:�<�
�w�}�#���6����	[�I�U���6�;�!�;�w�-�$���¹��^9��N��1��������}�BϺ�����O�
N��E��d�n�u�u�4�3����Y����g9��1��ڊ�&�
�u�u���8���&����|4�N�����u�|�o�u�g�m�F���s���P	��C��U����
�%�
�#�l����K����g"��x)��*�����}�u�8�3���Y���V��^�����u�:�&�4�#�<�(���	�֓�G��Q��F��������4���Y����\��XN�U��w�e�e�e�l�}�WϽ�����GF��h=�����&�2�
�&��}�W���&����p9��t:��U���1�"�!�u�~�g�W��I����l�N�����;�u�%���)�(���&����`2��{!��6�����u�`�3�*����P���W��^�N���u�6�;�!�9�}��������EU��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��h_��U���
���
��	�%���Y����G	�N�U��n�u�u�6�9�)����	����@��A_��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������ES��T��!�����
����_�������V�S��E��e�n�u�u�4�3����Y����\��h��G���o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�d�n�u�w�>�����ƭ�l��D��ߊ�e�o�����4���:����R��X����u�h�w�e�g��}���Y����G�������!�9�a�g�m��3���>����v%��eN��U���;�:�e�u�j��G��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���f�1�"�!�w�t�M���I����l�N�����;�u�%�6�9�)����O����g"��x)��*�����}�u�8�3���Y���W��UךU���:�&�4�!�6�����&����F��d:��9�������w�n��������\�_�E��u�u�6�;�#�3�W�������l
��h/��U���
���
��	�%���Y����G	�N�U��d�w�_�u�w�2����Ӈ��P	��C1��A���o������!���6�����Y��E���h�w�d�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�U�ԜY�Ư�]��Y�����;�!�9�a�f�g�$���5����l0��c!��]���:�;�:�e�w�`�U��H��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�f�1�"�#�}�^��Y����D��N�����!�;�u�%�4�3����M���5��h"��<������}�w�2����I����D��_�����u�:�&�4�#�<�(���
����9��N��1��������}�DϺ�����O�
N��D��n�u�u�6�9�)����	����@��AZ��U����
�����#���Q�ƨ�D��^��O���d�e�w�_�w�}��������C9��Y������o�����4���:����U��X����u�h�w�e�f�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�l�G���s���P	��C��U���6�;�!�9�b�o�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����lǻN�����9�4�
��1�0�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����]ǻN�����7�!�u�&��3��������G��PUךU���!�'�7�!�w�.�(�������	��V��&���8�o�&�2�6�}�������9F������4�
�<�
�$�,�$���¹��^9��N��1�����_�u�w�4��������T9��S1�U������n�w�}�����Ƽ�9��D�����
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h;�����1��e�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����,����_��~1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�;�4�1����I����E
��G��U����
���w�`�P���s���@��V��*ڊ�;�6�9�1��l��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�e� �&�4�2��(ށ����5��h"��<������}�b�9� ���Y���F�^�E��e�e�e�e�l�}�Wϭ�����C9��b ������
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G���
����W'��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�e��.����8����Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u����������lT��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�;�6�9�3��E���&����Z��^	��U���
���n�w�}�����Ƽ�9��D�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����R
��v'��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�֓�]��[��<���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�g��������� 9��h��*���&�2�o����0���s���@��V��*ڊ�;�6�9�1��n��������V�=��*����u�h�r�p�W�W���������h;�����1��a�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1�� ���4�0��
��/���*����|!��h8��!���}�`�1�"�#�}�^��Y����V��^�E��e�n�u�u�$�:����&ù��@��R
��*ފ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�e��.����8����R��[
�����o������M���I��ƹF��^	��ʥ�e� �&�4�2��(ځ�����\��c*��:���
�����h��������l�N�����u�
�
�;�4�1����L����TF��d:��9�������w�l�W������F��L�E��e�e�e�e�g��}���Y����R
��h^�����9�1��`�6���������\��c*��:���n�u�u�&�0�<�W���&����R
��v'��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u����������lP��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�G���
����W'��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�e� �&�6�8�6���&����_��Y1���������W�W���������h;�����1��c�4��1�(�������g"��x)��U��r�r�_�u�w�4����	�֓�]��[��<���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��D�����
�
�'�2�m��3���>����v%��eN��@ʱ�"�!�u�|�m�}�G��I����V��^�N���u�&�2�4�w��(�������r/��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�e� �&�4�2��(؁�	����l��PN�&������o�w�m�L���Yӕ��]��G1�� ���4�0��
��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*ڊ�;�6�9�1��e����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l3��T�����m�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u����������l^��G1�����0�u�u����>���D����l�N�����u�
�
�;�4�1����@����@��N��1��������}�F�������V�=N��U���;�9�%�e��.����8����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��E���&�4�0�����������@��N��1�����_�u�w�4����	�֓�]��[��<���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�G���
����W'��^�����2�o�����4���:����W��S�����|�_�u�u�>�3�Ϯ�I����P��S/��Dڊ�'�2�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��d��Uʦ�2�4�u�
��3��������9��h��*���&�2�o����0���s���@��V��*ڊ�;�6�9�1��l�(�������A��N��1�����o�u�g�f�W���
����_F��1�����0��
�d�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��E���&�4�0���l����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l3��T�����d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�m�"�������z9��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�9�>����0����Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u����������lW��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�e� �&�4�2��(�������W9��h��U����
���l�}�Wϭ�����C9��b ������
�g�4��1�(�������g"��x)��U��r�r�_�u�w�4����	�֓�]��[��<��
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lV��Y������d�
�'�0�g�$���5����l0��c!��]���1�"�!�u�~�g�W��I����V��^�E��u�u�&�2�6�}�(߁�����V��h_�����9�
�;�&�0�g�$���5����l�N�����u�
�
�;�4�1����H����l��h���������g�W��B�����Y����� �&�4�0���C���&����	F��s1��2������u�f�}�������9F������%�e� �&�6�8�6���M����TF��d:��9�������w�l�W������F��L�E��e�e�e�e�g��}���Y����R
��h^�����9�1��d��-��������TF��d:��9����_�u�u�>�3�Ϯ�I����P��S/��Dފ�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������r/��1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&����R
��v'��@���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�e��.����8����l��A�����<�u�u����>��Y����Z��[N��E���&�4�0���h��������V�=��*����u�h�r�p�W�W���������h,��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ѓ�lV��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�@���I����E
��G��U����
���w�`�P���s���@��V��*݊�
�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h,��*���2�o�����4���:����W��S�����|�o�u�e�g�m�G��I����D��N�����4�u�
�
����������@��N��1�����_�u�w�4����	�ѓ�lW��G1�����0�u�u����>���D����l�N�����u�
�
�
��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*݊�
�
�'�2�m��3���>����v%��eN��@ʱ�"�!�u�|�m�}�G��I����V��^�N���u�&�2�4�w��(���&����_��Y1���������W�W���������h,��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u���(܁�����\��c*��:���
�����h��������l�N�����u�
�
�
��/���*����|!��h8��!���}�`�1�"�#�}�^��Y����V��^�E��e�n�u�u�$�:����&Ĺ�� 9��h��*���&�2�o����0���s���@��V��*݊�
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u���(ہ����5��h"��<������}�b�9� ���Y���F�^�E��e�e�e�e�l�}�Wϭ�����C9��u1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��B���`�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(ځ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��7���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b��c�6���������\��c*��:���n�u�u�&�0�<�W���&����R��[
�����o������M���I��ƹF��^	��ʥ�b��b�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��7���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�`��@���&����Z��^	��U���
���n�w�}�����Ƽ�9�� 1��*���
�'�2�o���;���:���V�=N��U���;�9�%�b��e��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�b��m�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����;�ޓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��7���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�@���@����@��N��1��������}�F�������V�=N��U���;�9�%�b��d����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�w�_�w�}����Ӗ��l$��h�����<�
�<�u�w�	�(���0��ƹF��^	��ʥ�b��l�4��1�(�������g"��x)��U��r�r�_�u�w�4����	�ѓ�lW��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(؁�&�֓�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*���e�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���d�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��u1�*���2�o�����4���:����W��S�����|�o�u�e�g�m�G��I����D��N�����4�u�
�
��l��������l��T��!�����n�u�w�.����Y����q9��h�����%�0�u�u���8���Y���A��N�����4�u�
�
��o��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�b��d�
�%�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�M���I����V��^�E��n�u�u�&�0�<�W���&����l��A�����<�u�u����>��Y����Z��[N��B���d�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����l��D��Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�j�5��&����\��c*��:���
�����h��������\�^�E��e�e�e�e�g�f�W���
����_F�� 1��Dي�%�#�1�<��4�W���-����t/��=N��U���;�9�%�b��l�(�������A��N��1�����o�u�g�f�W���
����_F�� 1��Dފ�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��l$��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b��d��-��������TF��d:��9����_�u�u�>�3�Ϯ�N����9��h��*���2�o�����4��Y���9F������%�b��d��3����Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*݊�
�`�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�@���Hƹ��l��h�����o������}���Y����R
��hY��*���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�N���I����@��N��1��������}�D�������V�=N��U���;�9�%�l��m����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�@����l��A�����u�u��
���W��^����F�D�����
�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��D���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��z1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ʹ��9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����4�ԓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��8���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�N���J����@��N��1��������}�D�������V�=N��U���;�9�%�l��n����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�@����l��A�����u�u��
���W��^����F�D�����
�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��A���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��z1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ʹ��9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����4�ӓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��8���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�N���O����@��N��1��������}�D�������V�=N��U���;�9�%�l��k����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�@����l��A�����u�u��
���W��^����F�D�����
�
�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��B���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��z1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ʹ��9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����4�ޓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��8���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�N���@����@��N��1��������}�D�������V�=N��U���;�9�%�l��d����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�
�
�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�@����l��A�����u�u��
���W��^����F�D�����
�
�
�e�>�����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��L���d�
�'�2�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���Yӕ��]��G1��8��
�%�#�1�>�����Y����)��tUךU���<�;�9�%�n��F߁�	����l��PN�&������o�w�m�L���Yӕ��]��G1��8��
�;�&�2�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������l_��h_�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӗ��l+��1��*���
�;�&�2�m��3���>����F�D�����
�
�
�d�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l+��1��*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}�(ց�&�ԓ�C9��S1��*���u�u��
���L���Yӕ��]��G1��8��
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(ց�&�Փ�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�n��F܁����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�l��l�(�������]9��PN�&������_�w�}����Ӗ��l+��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�l��l�(���
���5��h"��<������}�f�9� ���Y����F�D�����
�
�
�a�'�8�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��P ��U���
�
�a�4��1�(���
���5��h"��<��u�u�&�2�6�}�(ց�&�ғ�C9��S1�����u��
���}�J���^���F��P ��U���
�
�`�<��4�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��8��
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��Dߊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�l��l�(�������A��N��1�����o�u�g�f�W���
����_F��1������
� �3�%�l�(���&����	F��s1��2������u�d�}�������9F������%�a��4�2��(�������9��P1�F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������z9��Q��*���g�'�2�c�a�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h=������7�3�0��h�E�������\��c*��:���
�����l��������l�N�����u�
�
�6�;�9�>�������R��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��h�����d�
�
�0��j�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��&���0��
� �1�/�Fہ�&����^��N��1��������}�D�������V�=N��U���;�9�%�a��<����&����V��1�����b�d�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�P��S/�����0�
�a�d��8�(��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������4�0���(����Hƹ��l��hY�U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������l��Q��Dފ�a�'�2�b�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h=������7�3�0��h�Fہ����� F��d:��9�������w�n�W������]ǻN�����9�%�a��6�8�6�������lW��D1����c�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����_��~1�����
�f�&�'�0�j�N��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���9�1��7�1�8�(���
����lQ��T��!�����
����_������\F��d��Uʦ�2�4�u�
��>����0����U��[��*���
�e�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z9��E1�����
�0�
�d�w�}�#���6����e#��x<��Aʱ�"�!�u�|�]�}�W�������A��B1�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����	F��s1��2������u�d�}�������9F������4�
�<�
�$�,�$���	ù��TT��D��U����
���l�}�Wϭ�����R��^	�����a�u�u����L���Yӕ��]��V�����%�!�;�%�g�4�G��*����|!��T��R��_�u�u�<�9�1��������l��h\�M��������4���Y����\��XN�N���u�&�2�4�w�-��������`2��G^�����3�8�a�o���;���:���F��P ��U���&�2�7�1�b�h�MϜ�6����l�N�����u�'�
� �o�m����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����g�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����&�2�
�&��}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��8�(�������CV��C_��U���
���u�j�z�P�ԜY�ƿ�T�������7�1�c�f�m��8���7���F��P ��U���!�:�1�
�"�e�A���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�%�&�2�2�4����H����lT��1��E���d�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��X��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���&����V��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(���A�ԓ�F��d:��9�������w�m��������l�N�����u�0�
�8�e�/���L����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�a�3��k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
�0�
�g�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1��܊� �m�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����g�b�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��Mڊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l��h\�E��������4���Y����\��XN�N���u�&�2�4�w�8�(���H����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�ށ�����Q�=��*����
����u�W������]ǻN�����9�&�9�!�'����K����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�f�%�:�E��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��&���
�:�
�:�'�l�(߁�����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������\��1�����'�2�g�e�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Z1��d;��:���&�3�
�e�a�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��^9��&����!�&�'�0�o�F���Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����%�f�3�
�g�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
�0�
�f�h�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���!�
�0�
�:�l�(���&����l��h��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����M����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����W��T��!�����
����_�������V�=N��U���;�9�4�
�2�����&����G��1����g�
�%�
�#�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Dߊ� �d�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��@���2�g�f�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��A��G�����9�!�%�`�%�:�E��&����Z��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�k����K����	F��s1��2������u�g�9� ���Y����F�D�����%�'�2�%�$�:��������l��h\�@���e�<�d�o���;���:����g)��^�����:�e�n�u�w�.����Y����G�� 1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��*��f�o�����4���:����V��X����n�u�u�&�0�<�W�������C��h��*���d�
�0�
�f�n�������5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�m�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���
�%�!�
�2����&����W��h��*���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}��������A��_�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�����	����@��C��L���2�g�c�
�'�����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������:�
�:�%�f��(���&����^��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��1�(���&����lW��1�����2�g�b�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƥ�l��u����
�
� �d�o��E��*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T�������,� �
�b�f�/���A����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʼ�
�<��'��2�(ځ�&¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�>���������C9��1�����g�m�u�u���8���&����|4�N�����u�|�_�u�w�4��������W��R��F���
�f�e�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��^	������
�%�
�#�l����K����g"��x)��N���u�&�2�4�w�-�������� ^�,��9���n�u�u�&�0�<�W�������G��hZ�����
�f�a�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��d�����
� �3�'�f��(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
�4�1��������A9��h_�����g�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�P��S/�����0�
�a�a�1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a��4�0����������9��P1�E���u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����r/��B����
�
� �d�c��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���9�1��7�1�8�(���A����lT��N�&���������W��Y����G	�UךU���<�;�9�%�c�����8����U ��h_��Dي� �d�b�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h=������7�3�0��i�F܁�����^�=��*����
����u�FϺ�����O��N�����4�u�
�
�4�1��������A9��h\�����a�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��V��4��� �3�'�d��l����K����	F��s1��2������u�d�}�������9F������%�a��4�2��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�P��S/�����0�
�a�g��8�(��A����g"��x)��*�����}�d�3�*����P���F��P ��U���
�6�9�1��?����&�ғ�9��h_�B���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��h�����d�
�a�'�0�o�D���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���4�0��
�"�;���&�ד�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������z9��Q��*���a�
�0�
�e�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hZ�����1��7�3�2��B�������U��N�&���������W��Y����G	�UךU���<�;�9�%�c�����8����U ��h_��D���2�g�a�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��V��4��� �3�'�d�����OĹ��\��c*��:���
�����l��������l�N�����u�
�
�6�;�9�>�������S��h��*��m�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����_��~1�����
�`�m�3��h�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������4�0���(����Hƹ��A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������l��Q��Dߊ�f�3�
�c�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��&���0��
� �1�/�Fځ�J����lT��N�&���������W��Y����G	�UךU���<�;�9�%�c�����8����U ��h_��Gۊ� �d�`�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h=������7�3�0��h�E؁����� 9��T��!�����
����_������\F��d��Uʦ�2�4�u�
��>����0����U��[��A���
�b�g�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��d�����
� �3�'�f��F���&����l��N��1��������}�D�������V�=N��U���;�9�<�
�>���������C��Q��G؊�a�o�����4���:����R��X����n�u�u�&�0�<�W���
����@��d:��Ҋ�&�
�u�u���8���B�����Y�����<�
�1�
�f�}�W���5����9F������2�%�3�
�d��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���m�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��hV�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_�������V�=N��U���;�9�:�
�8�9����Iǹ��\��c*��:���
�����}�������9F������;�"�0�
�"�e�O���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����0�d�3�
�f��D��*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T�������d�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��؊� �l�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V��[\�� ��g�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����V
��Q��Fފ�f�o�����4���:����W��S�����|�_�u�u�>�3�ϱ�&���� 9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}����ǹ��l_��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��1�(���@�֓� F��d:��9�������w�l�W������]ǻN�����9�;�"�0�o�;�(��&���5��h"��<������}�b�9� ���Y����F�D�����0��9�
�"�d�E���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����0�d�
� �n�e����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����d�
� �l�c�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��Y����
� �d�e��n�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��R�����3�
�e�m�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1��݊� �d�g�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��L���
�e�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��E���
�e�m�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��D���
�e�`�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��G���
�e�g�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����]��R�����c�
�f�o���;���:����g)��_����!�u�|�_�w�}����ӈ��`��1��*��e�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����Z9��E1�����
�
�g�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�
�:�1�
�"�l�Eف�K����g"��x)��*�����}�u�8�3���B�����Y�����0�d�
� �f�o�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V�����9�`�3�
�f�o����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��*���1�
� �d�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��X�����
� �d�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��@=��D܊� �d�a�
�d�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������d��B���
�d�c�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����\��X ��*���d�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�D5��V�� ��c�
�f�o���;���:����g)��_����!�u�|�_�w�}����ӈ��`��1��*��c�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����V
��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������_T��Q��D���%�u�u����>���<����N��
�����e�n�u�u�$�:��������U��B1�Eފ�f�o�����4���:����W��S�����|�_�u�u�>�3�ϰ�����9��h_�E���u�u��
���(���-���S��X����n�u�u�&�0�<�W���*����l ��\�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������U��\�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��[�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��X�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��X�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}�����֓�F9��Z��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���KĹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������l��Q��Dފ�
� �d�d��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hZ�����1��7�3�2��C�������_��N�&���������W��Y����G	�UךU���<�;�9�%�c�����8����U ��h_��B���
�f�c�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��d�����
� �3�'�f��G���&����l��N��1��������}�D�������V�=N��U���;�9�%�a��<����&����V��1�*���d�`�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lR��T�����7�3�0�
�c�l�(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
�4�1��������A9��h_�����f�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��V��4��� �3�'�d��e����J�ӓ� F��d:��9�������w�n�W������]ǻN�����9�%�a��6�8�6�������lW��W�� ��l�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l5��[��<���3�0�
�a�e����@ʹ��\��c*��:���
�����l��������l�N�����u�
�
�6�;�9�>�������R��1��*��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����`��R
��*���3�'�d�
�d�;�(��I����	F��s1��2������u�d�}�������9F������%�a��4�2��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�P��S/�����0�
�a�g��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����
�
�6�9�3���������lT��Q��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����&ǹ��R
��v'�� ���'�d�
�m�1��C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a��4�0����������_��B1�C؊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����_��~1�����
�a�f�
�"�l�Aց�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�6�9�1��?����&�ғ�9��h_�C���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��h�����d�
�g�3��i�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������4�0���(����Hǹ��l ��Z�*��o������!���6���F��@ ��U���_�u�u�<�9�1����*����W'��U�����a�f�
� �f�m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ފ�6�9�1��5�;����M����U��_�����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����r/��B����
�b�3�
�b�e����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���4�0��
�"�;���&�ޓ�F9��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������z9��Q��*���f�
� �d�d��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���9�1��7�1�8�(���Mù��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������l��Q��Dߊ�
� �d�c��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hZ�����1��7�3�2��B�������R��N�&���������W��Y����G	�UךU���<�;�9�%�c�����8����U ��h_��B���
�`�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��d�����
� �3�'�f��G���&����l��N��1��������}�D�������V�=N��U���;�9�%�a��<����&����V��1�*���d�e�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lR��T�����7�3�0�
�b�l�(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
�4�1��������A9��h_�����c�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��V��4��� �3�'�d��e����O�֓� F��d:��9�������w�n�W������]ǻN�����9�%�a��6�8�6�������lW��W�� ��f�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l5��[��<���3�0�
�`�e����Mǹ��\��c*��:���
�����l��������l�N�����u�
�
�6�;�9�>�������S��1��*��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����`��R
��*���3�'�d�
�d�;�(��L����	F��s1��2������u�d�}�������9F������%�a��4�2��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�P��S/�����0�
�`�g��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����
�
�6�9�3���������lT��Q��C���%�u�u����>���<����N��
�����e�n�u�u�$�:����&ǹ��R
��v'�� ���'�d�
�m�1��@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a��4�0����������_��B1�E݊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����_��~1�����
�`�f�
�"�l�Fہ�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�6�9�1��?����&�ӓ�9��h_�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��h�����d�
�g�3��j�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������4�0���(����Hƹ��l ��Y�*��o������!���6���F��@ ��U���_�u�u�<�9�1����*����W'��U�����`�f�
� �f�i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ފ�6�9�1��5�;����L����U�� [�����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����r/��B����
�b�3�
�`�n����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���4�0��
�"�;���&�ޓ�F9�� ^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������z9��Q��*���f�
� �d�`��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���9�1��7�1�8�(���Mù��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���A�ғ�VF��d:��9����_�u�u�>�3�Ͽ�&����@�=��*����
����u�W������]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����\��x!��4��u�u�&�2�6�}��������l_��T��:����n�u�u�$�:����	����l��hZ�Oʗ����_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����d�e�o����9�ԜY�ƿ�T�������7�1�d�l�m��8���7���F��P ��U���&�2�7�1�f�e�MϜ�6����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w�-��������F��u!��0���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:����	����l��hX�Oʗ����_�w�}����Ӈ��@��U
��B���u����l�}�Wϭ�����R��^	�����c�o�����}���Y����R
��G1�����1�l�u�u���6��Y����Z��[N��*���
�1�
�e�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��l�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&���� V��N��:����_�u�u�>�3�Ͽ�&����Q��_�Oʗ����_�w�}����Ӈ��@��U
��F���o�����W�W���������D�����f�a�o����9�ԜY�ƿ�T�������7�1�f�f�m��8���7���F��P ��U���&�2�7�1�d�o�MϜ�6����l�N�����u�%�&�2�5�9�E��CӤ��#��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���
����W��]��U�����n�u�w�.����Y����Z��S
��C���u����l�}�Wϭ�����R��^	�����b�u�u����L���Yӕ��]��V�����1�
�m�u�w��;���B�����Y�����<�
�1�
�o�}�W���5����9F������4�
�<�
�3��N���Y����v'��=N��U���;�9�4�
�>�����O����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�L������]�}�W�������C9��P1����m�o�����}���Y����R
��G1�����1�a�b�o���2���s���@��V�����2�7�1�a�a�g�5���<����F�D�����%�&�2�7�3�n�G��;����r(��N�����4�u�%�&�0�?���@����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lU��T��:����n�u�u�$�:����	����l��hZ�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�g�u�u���6��Y����Z��[N��*���
�1�
�f�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��i�W���6����}]ǑN�����:�0�!�8�e�l�3۟�&ù��F
�� ��Fػ�
�g�d�8�/�9�ϗ�s���T��E��]���u�u�u��w�}�9���<��ƹF�N�� �����u�u���2��Y���F��^ ��"����o�����}���Y���W��h9��!���u����l�}�W���Yӂ��G9��s:��Oʜ����|�]�}�W�����ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}����Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����u�u� �u���8���&����|4�_�����:�e�u�n�w�}��������]��dװU���6�8�:�0�#�0�E��=ǧ��9��C��*���
�g�g��]�}�W�������l�N��Uʜ�u�u����f�W���Y����f+��c/��U������n�w�}�W�������d/��N�<�����_�u�w�}�W�������g.�'��0���u�n�u�u�'�/�W�ԜY���F��\N�<����
���l�}�W���YӔ��V�'��&������_�w�}�W������/��d:��9�������w�n�W������]ǻN��U���0�o��u���8���B���F�
����������4���:����U��S�����|�|�_�u�w�3�W���	����G]Ǒ=d�����u�u�3�e�1�(�(���
����@9��h_�����&�
�e�o�4�0����Ӌ��W��/��E��� �
�g�&�d�3�(���H����l��=N��U���0�<�u�4�w�W�W���Y�ƅ�[�BךU���u�u� �
���W���H���F�N��ڊ���u�k�d�q�W���Y����Z��`'��=��u�g�_�u�w�}�W�������g.�	N�\���u�%�'�u�6�}�}���Y���W��S����3�
�f�
�g�W�W���Y�ƨ�]W�	N�����
�f�
�d�]�}�W���Y����[�P�����f�
�g�n�]�}�W���&����U����G��� �u�u�:�'�3����;����wR��h^�����%�f�&�f��W�W�������PF��GN��U���u�u��u�i�l�}���Y���}3��d:��0��u�y�u�u�w�}����&����{F�]����u�u�u�:�#�
�3���D����l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N����h�u�'�
�"�e�C���U���F���H���'�
� �m�c�>�[���Y�����CN��U���
� �m�a�'�t�}�Զs���K�C�����0�!�&�4�2�u����&����	��C�����0�8�6�<�2�}�Z���YӇ��p5��D�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�_�u�w�}�W���Y���F�V��&���8�i�u�%�����Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�4�
�2���������l�������%�:�0�&�w�p�W�������T9��^��*���
�!�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W�������C��Y1��E���e�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Yۇ��@��U
��D��|�!�0�u�w�}�W���Y���F�N��U���%�'�2�%�>�8�(���&����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���O�Ƹ�V�N��U���u�u�u�u�w�}�W�������T9��^��*���
�!�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w�-����	����]9��1��Dʴ�&�2�u�'�4�.�Y��s���R��R	�����;�%�e�<�f�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӇ��A��G�����%�
�!�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N�����-�!�:�1��8�(��A����C9��Y�����e�u�;�u�6�����&����P9��
N��*���
�&�$���-�(���J����lR�N�����u�u�u�u�w�}�W���Y����C9��P1�����
�%�
�!�w�`��������_	��T1����u�u�u�u�w�}�W������N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lW������4�1�;�!�6��������� O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����&�2�
�&��t�������V��T��D���2�g�f�u�w�-��������lV�G�����u�u�u�u�w�}�W���Y�����E�����0�
�%�
�#�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��Y������e�4�
�;���������]F��X�����x�u�u�%�g���������9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G���
����W'��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��CV�����|�u�=�;�]�}�W���Y���F�N��U���%�e� �&�6�8�6���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR�����ߊu�u�u�u�w�}�W���Y���F��1�����0��
�
�'�+���������h;�����1��e�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�;�6�9�3��G����ƭ�@�������{�x�_�u�w��(�������r/��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g���������9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�
��3��������l��A��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(������O��_�����u�u�u�u�w�}�W���Y����f��V��4���
�'�2�i�w��(�������r/��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�e� �$�<����&�֓�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u����������lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�e� �&�4�2��(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����U�����ߊu�u�u�u�w�}�W���Y���F��1�����0��
�e�6��������F��1�����0��
�e�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�;�6�;�9�>��&������^	�����0�&�u�x�w�}����,����_��~1�*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G���
����W'��^�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�e� �$�<����&�֓�C9��SG��U���;�_�u�u�w�}�W���Y���F��1�����0��
�e�'�8�W��	�֓�]��[��<��n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����0��
�d�6���������@��YN�����&�u�x�u�w�-�G���
����W'��_�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��@��R
��*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N��U���u�u�u�%�g���������W��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��Uʥ�e� �&�4�2��(�������W9��R	��Hʥ�e� �&�4�2��(�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������lW��G��U���<�;�%�:�2�.�W��Y����lV��Y������d�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l3��T�����d�
�'�2�k�}��������EW��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�G���
����W'��_�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e� �&�4�2��(���	����[��h^�����9�1��d�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(�������W9��R	�����;�%�:�0�$�}�Z���YӖ��l3��T�����d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����0��
�g�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�u�u�u�w�}�WϮ�I����P��S/��D؊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�d�l�w�5��ԜY���F�N��U���u�u�u�%�g���������T��G1�����0�u�h�%�g���������T��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���%�0�u�&�>�3�������KǻN��*ڊ�;�6�9�1��l�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���6�9�1��f�����E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l3��T�����d�
�%�#�3�t�W������F�N��U���u�u�u�%�g���������T��E��I���
�
�;�6�;�9�>��B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g���������U��G1�����0�u�&�<�9�-����
���9F���*���6�9�1��f���������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�e� �&�4�2��(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�}�W���Y�����h;�����1��d�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�F��Y����l�N��U���u�u�u�u�w�}�WϮ�I����P��S/��Dي�%�#�1�%�2�}�JϮ�I����P��S/��Dي�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����0��
�f�'�8�W�������A	��D�X�ߊu�u�
�
�9�>����0����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�;�4�1����H����V�
N��*���&�
�#�c�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���6�9�1��f��������G��d��U���u�u�u�u�w�}�WϮ�I����P��S/��Dي�'�2�i�u����������lW��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�I����P��S/��Dފ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�;�4�1����Hǹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g���������R��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��Q��@���!�0�u�u�w�}�W���Y���F�N��U���
�;�6�9�3��Fہ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������Q�C��U���u�u�u�u�w�}�W���Y�����h;�����1��d�
�'�+���������h;�����1��d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(���	����R��P �����&�{�x�_�w�}�(߁�����V��h_�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������r/��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�;�4�1����Hǹ��l��G�����u�u�u�u�w�}�W���Y�����h;�����1��d�
�%�:�K���&ù��@��R
��*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h;�����1��d�
�'�+�����ƭ�@�������{�x�_�u�w��(�������r/��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�I����P��S/��Dߊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
��3��������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��B���!�0�u�u�w�}�W���Y���F�N��U���
�;�6�9�3��Fځ�	����l��PN�U���
�;�6�9�3��Fځ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g���������S��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�`�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����f��V��4���`�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������r/��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�;�6�9�3��Fځ����F��1�����0��
�`�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�;�6�9�3��F���&����C�������%�:�0�&�w�p�W���	�֓�]��[��<���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��Y������d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��U���u�u�u�u�w�-�G���
����W'��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����e�u�=�;�]�}�W���Y���F�N��U���%�e� �&�6�8�6���&����_��E��I���
�
�;�6�;�9�>�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������lW��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�]��[��<���%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������lW��G1�����u�=�;�_�w�}�W���Y���F�N��E���&�4�0�������E�Ƽ�9��D�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
��-����	����R��P �����&�{�x�_�w�}�(߁�����V��h\�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��@��R
��*؊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
��3��������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ڊ�;�6�9�1��o��������V�
N��E���&�4�0����������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e� �$�<����&����V��D��ʥ�:�0�&�u�z�}�WϮ�I����P��S/��G���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(߁�����V��h\�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�e� �$�<����&����l��G�����u�u�u�u�w�}�W���Y�����h;�����1��g�%�2�}�JϮ�I����P��S/��G�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��Y������f�4�
�;���������]F��X�����x�u�u�%�g��������� 9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G���
����W'��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��CV�����|�u�=�;�]�}�W���Y���F�N��U���%�e� �&�6�8�6���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lP�����ߊu�u�u�u�w�}�W���Y���F��1�����0��
�
�'�+���������h;�����1��f�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�;�6�9�3��D����ƭ�@�������{�x�_�u�w��(�������r/��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g��������� 9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�;�6�9�3��D���&����O��_�����u�u�u�u�w�}�W���Y����f��V��4���
�'�2�i�w��(�������r/��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*ފ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�;�4�1����M����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��3��������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ڊ�;�6�9�1��i��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l3��T�����a�4�
�9��/���Y����f��V��4���
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
��/�Ͽ�
����C��R��U���u�u�%�e��.����8����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�;�4�1����M����TF������!�9�d�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1�� ���4�0��
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����,����_��~1�����u�h�%�e��.����8����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�G���
����W'��1��*���
�'�2�4�$�:�W�������K��N����� �&�4�0���(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e� �&�6�8�6���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���A����lS����ߊu�u�u�u�w�}�W���Y���F��1�����0��
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�O�������9F�N��U���u�u�u�u�w�}�W���&����R
��v'��*���#�1�%�0�w�`����,����_��~1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��Y������`�%�0�w�.����	����@�CךU���
�
�;�6�;�9�>���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N����� �&�4�0���(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��Y������`�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u����������lS��E��I���
�
�;�6�;�9�>��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��3��������l��A�����u�&�<�;�'�2����Y��ƹF��h^�����9�1��c�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�;�6�9�1��k��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l3��T�����c�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�b�}����s���F�N��U���u�u�u�u�'�m�"�������z9��V�����'�2�i�u����������lP��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*܊�'�2�4�&�0�}����
���l�N��E���&�4�0�����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^�����9�1��c�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ù��@��R
��*܊�%�#�1�|�w�5��ԜY���F�N��U���u�%�e� �$�<����&Ź��V�
N��E���&�4�0���f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�e� �&�6�8�6���&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����0��
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�m�1�0�B�������9F�N��U���u�u�u�u�w�}�W���&����R
��v'��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�a�u�?�3�}���Y���F�N��U���u�u�%�e��.����8����R��[
�����i�u�
�
�9�>����0�ѓ�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����V��hY�����4�&�2�u�%�>���T���F��1�����0��
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��Y������b�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(߁�����V��hY�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e� �&�4�2��(؁����F��1�����0��
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C���� �&�4�0���(�������A��V�����'�6�&�{�z�W�W���&ù��@��R
��*Ҋ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��D�����
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�b�t����Y���F�N��U���u�u�u�u�w��(�������r/��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����f�u�=�;�]�}�W���Y���F�N��U���%�e� �&�6�8�6���&����_��E��I���
�
�;�6�;�9�>�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������l^��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�]��[��<���%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������l^��G1�����u�=�;�_�w�}�W���Y���F�N��E���&�4�0�������E�Ƽ�9��D�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
��-����	����R��P �����&�{�x�_�w�}�(߁�����V��hW�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��@��R
��*ӊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
��3��������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�G���=�;�_�u�w�}�W���Y���F�N����� �&�4�0���(�������A��S��*ڊ�;�6�9�1��d������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�9�>����0�ߓ�A��V�����'�6�&�{�z�W�W���&ù��@��R
��*ӊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����,����_��~1�����u�h�4�
�8�.�(���O����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�9�>����0�ߓ�C9��SG��U���;�_�u�u�w�}�W���Y���F��1�����0��
�
�%�:�K���&ù��@��R
��*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��u1�����9�
�'�2�6�.��������@H�d��Uʥ�b��e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���m�3�8�`�~�)����Y���F�N��U���u�u�u�u���(߁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������Q�C��U���u�u�u�u�w�}�W���Y�����h,��*���#�1�%�0�w�`����;�֓�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(؁�&ù��V��D��ʥ�:�0�&�u�z�}�WϮ�N����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b��g�-����DӇ��P	��C1��D܊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����q9��V�����|�!�0�u�w�}�W���Y���F�N��*݊�
�
�'�2�k�}�(؁�&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�5��&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��^�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��V��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��Q��@���!�0�u�u�w�}�W���Y���F�N��U���
�
�e�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��G�������9F�N��U���u�u�u�u�w�}�W���&����l��A�����u�h�%�b��l�(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��l�(���Ӈ��Z��G�����u�x�u�u�'�j�5��&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�e�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����l��A��\���=�;�_�u�w�}�W���Y���F�G1��7��
�'�2�i�w��(���I���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(�������W9��R	�����;�%�:�0�$�}�Z���YӖ��l$��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N����9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����G^��D��\���=�;�_�u�w�}�W���Y���F�N������d�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�A������F�N��U���u�u�u�u�w�}����;����R��[
�����i�u�
�
��l������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��l����Y����T��E�����x�_�u�u���(���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������d�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����;����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hY��*���%�0�u�h�'�j�5��B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`��F݁�	����l��PN�����u�'�6�&�y�p�}���Y����q9��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�
�g�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��o�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&�ԓ�C9��S1�����h�%�b��f��������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�b��f���������]F��X�����x�u�u�%�`��F݁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�g�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�&�ԓ�C9��SG��U���;�_�u�u�w�}�W���Y���F�� 1��D؊�'�2�i�u���(��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
���D���&����C�������%�:�0�&�w�p�W���	�ѓ�lW��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����;����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����l ��h[��U���;�_�u�u�w�}�W���Y���F�N��B���d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�d�i�W������F�N��U���u�u�u�u�w�-�@���H����l��h����u�
�
�
�d�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
�d�-����
������T��[���_�u�u�
���D�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���d�
�'�2�k�}��������EW��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@���H����l��G�����u�u�u�u�w�}�W���Y�����h,��F���0�u�h�%�`��F��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��l�(�������A��V�����'�6�&�{�z�W�W���&Ĺ��R��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�&�ғ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�W���Y���F���*���a�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�c�t����Y���F�N��U���u�u�u�u�w��(���M����E
��G��U��%�b��d��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��d��/�Ͽ�
����C��R��U���u�u�%�b��l�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���a�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(���M����E
��G�����_�u�u�u�w�}�W���Y���C9��u1�*���2�i�u�
���C�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��h��������V��D��ʥ�:�0�&�u�z�}�WϮ�N����9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@���Hƹ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����_�u�u�u�w�}�W���Y���F�G1��7��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�f�e�}����s���F�N��U���u�u�u�u�'�j�5��&����_��E��I���
�
�
�`�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�`�'�8�W�������A	��D�X�ߊu�u�
�
��h����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��7��
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�5��&����_�N�����u�u�u�u�w�}�W���Y����lQ��h_�����u�h�%�b��l�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�b��f�<�(���&������^	�����0�&�u�x�w�}����;�ד�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(ށ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�}�W���Y���C9��u1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�g�|�!�2�}�W���Y���F�N��U���u�u�
�
����������TF���*���
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��7���%�0�u�&�>�3�������KǻN��*݊�
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�lW��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�b��d�4��1�^�������9F�N��U���u�u�u�u�w��(���&����Z�G1��7��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h,��*���#�1�%�0�w�.����	����@�CךU���
�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���g�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N��U���u�u�u�u�'�j�5�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����U�����ߊu�u�u�u�w�}�W���Y���F�� 1��G���
�9�
�'�0�a�W���&����R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����;�ԓ�A��V�����'�6�&�{�z�W�W���&Ĺ��9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l$��h�����|�u�=�;�]�}�W���Y���F�N������g�%�0�w�`����;����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�N����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�e�i�W������F�N��U���u�u�u�u�w�-�@���J����E
��G��U��%�b��f�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�%�:�����Ƽ�\��D@��X���u�%�b��d�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1��F���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������F��R ��U���u�u�u�u�w�}�W���	�ѓ�lU��E��I���
�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����a�4�
�;���������]F��X�����x�u�u�%�`��C���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�o�;���PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��@���!�0�u�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����lQ��hZ�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��1�����&�<�;�%�8�8����T�����h,��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@���M����TF������!�9�d�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��7���4�
�9�|�~�)����Y���F�N��U���u�u�
�
������E�Ƽ�9��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�lS��G1�����0�u�&�<�9�-����
���9F���*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��u1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F�N��U���u�%�b��b�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����O����[��=N��U���u�u�u�u�w�}�W���Y����q9��V�����'�2�i�u���(ځ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`��B����ƭ�@�������{�x�_�u�w��(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����;�ӓ�C9��SG��U���;�_�u�u�w�}�W���Y���F�� 1��@���0�u�h�%�`��B�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
����������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�5�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�}�W���Y�����h,��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�g�d�u�?�3�}���Y���F�N��U���u�u�%�b��k��������V�
N��B���c�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�'�2�4�$�:�W�������K��N������c�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����q9��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�@���O����TF���*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1��B���
�9�
�'�0�<����Y����V��C�U���%�b��b�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�b�t����Y���F�N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lT��N�����u�u�u�u�w�}�W���Y���F��hY��*݊�%�#�1�%�2�}�JϮ�N����l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����C�������%�:�0�&�w�p�W���	�ѓ�lQ��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b��j����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9�� 1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�
�'�0�a�W���&����9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@���A����E
��G��U���<�;�%�:�2�.�W��Y����lQ��hV�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����G^��D��\���=�;�_�u�w�}�W���Y���F�N������m�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��e�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&˹��l��h����u�
�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��m�'�8�W�������A	��D�X�ߊu�u�
�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hY��*Ҋ�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`��O���&����O��_�����u�u�u�u�w�}�W���Y����q9��G��U��%�b��m�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�
�%�!�9����Y����T��E�����x�_�u�u���(ց�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b��n�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�l_��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��G��u�=�;�_�w�}�W���Y���F�N��Uʥ�b��l�4��1�(������C9��u1�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��hW�����4�&�2�u�%�>���T���F�� 1��L���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�&ʹ��V�
N��*���&�
�#�c�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�}����s���F�N��U���u�u�%�b��d����Y����lQ��hW�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����~9��V�����'�2�4�&�0�}����
���l�N��L���e�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��M���8�`�|�!�2�}�W���Y���F�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����J���G��d��U���u�u�u�u�w�}�W���YӖ��l+��h�����%�0�u�h�'�d�:�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(߁�����@��YN�����&�u�x�u�w�-�N���I����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�l��e�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hW��*ڊ�'�2�i�u���(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�l��l�(�������A��V�����'�6�&�{�z�W�W���&ʹ��V��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ց�&�֓�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�W���Y���F���*���e�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�b�t����Y���F�N��U���u�u�u�u�w��(���I����E
��G��U��%�l��d��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�l��d��/�Ͽ�
����C��R��U���u�u�%�l��l�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���e�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(���I����E
��G�����_�u�u�u�w�}�W���Y���C9��z1�*���2�i�u�
���G�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��l��������V��D��ʥ�:�0�&�u�z�}�WϮ�@����9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�N���H¹��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����_�u�u�u�w�}�W���Y���F�G1��8��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�a�g�}����s���F�N��U���u�u�u�u�'�d�:��&����_��E��I���
�
�
�d�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�d�'�8�W�������A	��D�X�ߊu�u�
�
��l����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��8��
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:��&����_�N�����u�u�u�u�w�}�W���Y����l_��h_�����u�h�%�l��l�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l��f���������TF��D��U���6�&�{�x�]�}�W���&����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���K����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9��N�����u�u�u�u�w�}�W���Y���F��hW��*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�c�~�)����Y���F�N��U���u�u�u�u���(�������W9��R	��Hʥ�l��d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�l��d�
�%�:�����Ƽ�\��D@��X���u�%�l��f���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hW��*���%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���(�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��\�����i�u�
�
��o�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
�d�<�(���&������^	�����0�&�u�x�w�}����4����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�d�:��&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���A����lS����ߊu�u�u�u�w�}�W���Y���F��1��Dي�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�a�m�w�5��ԜY���F�N��U���u�u�u�%�n��F܁�	����l��PN�U���
�
�f�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�f�%�2�}����Ӗ��P��N����u�
�
�
�d�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1��Dي�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�n��F܁�	����O�C��U���u�u�u�u�w�}�W���YӖ��l+��1�����h�%�l��f�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�l��d��-����	����R��P �����&�{�x�_�w�}�(ց�&�ғ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�}�W���Y�����h#��A���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�}�W���YӃ��Z �V�����1�
�m�|�#�8�W���Y���F�N��U���u�u�u�
���C���&����C��R������d�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����d�
�'�0�<����Y����V��C�U���%�l��d��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h#��A���0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���C���&����O��_�����u�u�u�u�w�}�W���Y����~9��h����u�
�
�
�c�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�`�6���������@��YN�����&�u�x�u�w�-�N���Hƹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�n��Fځ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�}�W���Y���C9��z1�*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�a�c�u�?�3�}���Y���F�N��U���u�u�%�l��l�(�������A��S��*ӊ�
�`�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ӊ�
�`�%�0�w�.����	����@�CךU���
�
�
�`�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��z1�*���2�i�u�%�4�3����J����9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�l��l�(������F��R ��U���u�u�u�u�w�}�W���	�ߓ�lW��G��U��%�l��d�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�l��d�4��1�(���Ӈ��Z��G�����u�x�u�u�'�d�:�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�}�'�>��������lW������6�0�
��$�e����L����[��=N��U���u�u�u�u�w�}�W���Y����~9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�
�'�+���������h#��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��z1�����u�&�<�;�'�2����Y��ƹF��hW��*ۊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����4�ד�A��S�����;�!�9�f��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��L���d�4�
�9�~�t����Y���F�N��U���u�u�u�
���(������C9��z1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l+��h�����%�0�u�&�>�3�������KǻN��*ӊ�
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1��G���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:��Ҋ�&�
�|�u�?�3�}���Y���F�N��U���u�u�%�l��o��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�
9��1��*���
�'�2�i�w��(���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�:���	����R��P �����&�{�x�_�w�}�(ց�&����V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�@����l��A��\���=�;�_�u�w�}�W���Y���F�G1��8���%�0�u�h�'�d�:��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
���(�������A��V�����'�6�&�{�z�W�W���&ʹ�� 9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�N���J����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9��N�����u�u�u�u�w�}�W���Y���F��hW��*ي�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�f�m�w�5��ԜY���F�N��U���u�u�u�%�n��D���&����C��R������f�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ӊ�
�
�'�2�6�.��������@H�d��Uʥ�l��f�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�
9��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����4�Փ�A��S��*ӊ�
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��8���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�l��c�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�m�3�:�h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ց�&ǹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��Y�����u�u�u�u�w�}�W���Y���F���*���
�%�#�1�'�8�W��	�ߓ�lR��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ʹ��9��R	�����;�%�:�0�$�}�Z���YӖ��l+��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�n��C��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��z1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�
�%�:�K���&ʹ��]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����4�ӓ�C9��S1�����&�<�;�%�8�8����T�����h#��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����~9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�l��`�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��G�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�
�
���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�l��b�-����
������T��[���_�u�u�
���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��1�����h�%�l��b�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l��k��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l+��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����`�u�=�;�]�}�W���Y���F�N��U���%�l��c�6��������F��1��C���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h#��*���2�4�&�2�w�/����W���F�G1��8���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ӊ�
�
�%�#�3�t�W������F�N��U���u�u�u�%�n��A��������h#��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�
9�� 1��*���
�'�2�4�$�:�W�������K��N������b�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hW��*݊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
���(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����l_��hY�����1�%�0�u�j�-�N���N����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���&������^	�����0�&�u�x�w�}����4�ѓ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�l��b�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ʹ��9��h��\���!�0�u�u�w�}�W���Y���F���*���
�'�2�i�w��(���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�n��O���&����C�������%�:�0�&�w�p�W���	�ߓ�l^��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ց�&˹��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����_�u�u�u�w�}�W���Y���F�G1��8���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�f�~�)����Y���F�N��U���u�u�u�u���(ׁ�	����l��PN�U���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����m�%�0�w�.����	����@�CךU���
�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����l_��hV�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�l��o�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����C��R������m�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�l��l�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���u�u�u�u�w�}����4�ߓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��Z�U���;�_�u�u�w�}�W���Y���F�N��L���l�4�
�9��/���Y����~9��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�l_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(ց����F��h�����#�g�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h#��*���#�1�|�u�?�3�}���Y���F�N��U���%�l��l�'�8�W��	�ߓ�l_��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W�������A9��X��*���
�d�u�&�>�3�������KǻN��9���
�:�
�:�'�h����A�ޓ�@��Y1�����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�;�_���
����W��^�����u�u�u�u�w�}�W���Y�����[�����:�%�`�'�0�e�O��Y����Z9��E1�����
�
�
�0��l�O�ԜY���F�N��Uʰ�&�3�}�%�$�:����O���G��d��U���u�u�u�u�w�}�WϷ�&����\��X��@���2�m�m�i�w�-��������lV��N��U���u�u�u�u�2�9���Y���F�N�����3�u�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ڊ�!�e�3�8�f�t�W������F�N��U���u�%�'�2�'�.��������WW��R	��E���%�e�<�d�k�}��������A��^�N���u�u�u�u�w�}�WϿ�&����C��P1�����%�f�'�2�e�l�(���&����[��R����
�0�
�d�b�W�W���Y���F�N��*���
�%�!�
�2����&����W��h��*���u�h�&�9�#�-�C�������]ǻN��U���u�u�u�u�'�/����
����V
��Z�*���
�d�c�%�g�4�F��Y����G��1����f�n�u�u�w�}�W���Y����C9��P1�����&�9�!�%�a�/���Mƹ��9��N�U���
�8�d�
�2��F��s���F�N��U���4�
�0�
�'�)�(���&����9��P1�@ي�%�
�!�u�j�.����	�ѓ�V��[����u�u�u�u�w�}�W�������C��h��*���d�
�0�
�f�m�������F��[1�����'�2�g�c�l�}�W���Y���F������%�&�2�&�;�)��������P��G����i�u�0�
�:�l�(���&����l�N��U���u�u�u�0�>�>��������U��S�����:�1�
� �o�k���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��E���2�
�&�
�~�<����	����@��A_��U���-�!�:�1��(�O���	�����Yd��U���u�u�u�u�w�;�(���?����\	��Z��*���
�0�
�d�b�a�W�������A9��X��A���%�<�3�
�g�d���Y���F�N��U����9�
�:��2���&¹��Z9��P1�B���h�3�
�!��/�;���&�ғ�l��h��D��
�f�_�u�w�}�W���Y���Z1��d;��:���d�
�
�0��l�D��Y����`3��x��D݊�
� �d�m��o�}���Y���F�N��������!�$�/���H�����O=�����
�
� �d�a��E�ԜY���F�N��Uʦ�9�!�%�f�%�:�E��Y����V
��Z�*���d�b�
�g�]�}�W���Y���F�D�����a�'�2�g�e�}�Jϭ�����R��B1�Mފ�g�_�u�u�w�}�W���Y�ƿ�_9��G_�����g�f�u�h�$�1����L����V��h����u�u�u�u�w�}�W���&����9��P1�A���h�&�9�!�'�k����I�Г�]ǻN��U���u�u�u�u�2����&����W��R�����!�%�b�3��l�E���B���F�N��U���u�0�
�8�f�����H���F��[1�����3�
�d�m�'�f�W���Y���F�N�����8�d�
�0��l�A��Y����G��1��*��a�%�n�u�w�}�W���Y�����h��D���2�g�m�u�j�.����	¹��l^��h����u�u�u�u�w�}�W���&����l��h\�F��u�0�
�8�e�;�(��&����F�N��U���u�u�&�9�#�-�(���&����Z�D�����
� �m�g�'�f�W���Y���F�N�����8�a�'�2�e�k�W��
����^��Q��CҊ�g�_�u�u�w�}�W���Y�ƿ�_9��GX�����e�g�i�u�2���������9��d��U���u�u�u�u�w�.����	˹��T9��^��Hʦ�9�!�%�
�"�e�G���B���F�N��U���u�0�
�8��8�(��K���@��C�����`�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�'�0�-����&����Z����U´�
�:�&�
�8�4�(���Y����Z��D��&���%�
�!�e�1�0�F�������C9��Y�����e�h�0�<�4�3�F���&����CT�N���ߊu�u�u�u�w�}�W���5����u	��{��*ߊ�
�
�0�
�f�e�K���5����u	��{��*ߊ�
�
� �d�n��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������G��G����u�;�u�4��2��������F�V�����&�$��
�'���������F��SN�����;�!�9�d�g�`��������@��R�����d�'�2�g�d��߁������Yd��U���u�u�u�u�w�-�C�������z9��Q��*���&�'�2�b�a�a�W���&����V��h�����d�
�a�'�0�o�D��Y���F�N��U���
�
�6�9�3���������l��R	��B���h�%�a��6�8�6�������lW��Z�� ��a�
�f�_�w�}�W���Y���F��1������
� �3�%�l�(�������V�
N��A���4�0��
�"�;���&�ѓ�V��\����u�u�u�u�w�}�W���&����V��h�����d�
�c�'�0�j�C��Y����`��R
��*���3�'�d�
�f�/���K��ƹF�N��U���u�u�
�
�4�1��������A9��h\�����f�u�h�%�c�����8����U ��h_��A���2�g�e�n�w�}�W���Y���F��hZ�����1��7�3�2��C�������T�
N��A���4�0��
�"�;���&˹��T9��]�U���u�u�u�u�w�}����*����W'��U�����a�l�'�2�a�e�K���&ǹ��R
��v'�� ���'�d�
�f�%�:�E��B���F�N��U���u�
�
�6�;�9�>�������R��R	��D���h�%�a��6�8�6�������lW��1����e�n�u�u�w�}�W���Y����lR��T�����7�3�0�
�c�.����N���F��1������
� �3�%�l�(�������U��=N��U���u�u�u�u�w��(�������l��Q��Dߊ�a�'�2�b�d�a�W���&����V��h�����d�
�b�3��k�D���B���F�N��U���u�
�
�6�;�9�>�������S��1����b�i�u�
��>����0����U��[��D���
�c�d�%�l�}�W���Y���F���*���9�1��7�1�8�(���K����lP��R������4�0���(����Hƹ��A��\�N���u�u�u�u�w�}�WϮ�M����_��~1�����
�`�`�'�0�k�B��Y����`��R
��*���3�'�d�
��8�(��J���F�N��U���u�%�a��6�8�6�������lW��1����d�i�u�
��>����0����U��[��F���2�g�`�n�w�}�W���Y���F��hZ�����1��7�3�2��B�������Z�G1��&���0��
� �1�/�Fځ�&����T��d��U���u�u�u�u�w�-�C�������z9��Q��*���&�'�2�m�b�a�W���&����V��h�����d�
�d�3��j�F���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����C��R ��ڊ�!�|�4�1��%����¹��T9��V��U���6�;�!�9�f�m�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��P]�����|�|�!�0�]�}�W���Y���F�G1��&���0��
� �1�/�Fہ�J����lT��N�U���
�6�9�1��?����&�ғ� 9��h_�D���n�u�u�u�w�}�W���YӖ��l5��[��<���3�0�
�a�f�/���I�����h=������7�3�0��i�F���&����l��=N��U���u�u�u�u�w��(�������l��Q��Dފ�
�0�
�g�o�a�W���&����V��h�����d�
�
� �f�o�(��s���F�N��U���%�a��4�2��(�������9��E��G��u�h�%�a��<����&����V��1�����f�f�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۃ��G��S_�����e�m�h�4��2����¹����F��*���&�
�:�<��}�W���
����@��d:��ڊ�!�e�3�8�f�}��������]��[����h�4�
�0��-����	�֓�GW�N���ߊu�u�u�u�w�}�W���&ǹ��R
��v'�� ���'�d�
�d�%�:�E��Y����lR��T�����7�3�0�
�c�o�(���H����CU��N��U���u�u�u�u�'�i�$�������Q��R��A��
�0�
�g�o�a�W���&����V��h�����d�
�b�3��i�O���B���F�N��U���u�
�
�6�;�9�>�������R��1����f�u�h�%�c�����8����U ��h_��Fފ� �d�l�
�d�W�W���Y���F�N��A���4�0��
�"�;���&�ד�V��]�I���
�
�6�9�3���������lR��Q��@���%�n�u�u�w�}�W���Y����lR��T�����7�3�0�
�b�l�(���&����Z�G1��&���0��
� �1�/�Fځ�J����P��h����u�u�u�u�w�}�W���&����V��h�����d�
�
�0��o�D��Y����`��R
��*���3�'�d�
��(�F��&����F�N��U���u�u�%�a��<����&����V��1�����g�a�u�h�'�i�$�������Q��R��@���3�
�`�b�'�f�W���Y���F�N��*ފ�6�9�1��5�;����L�ޓ�V��[�I���
�
�6�9�3���������l^��B1�MҊ�f�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���	ù��TT��D��\ʴ�1�}�-�!�8�9�(���&����[��G1�����9�d�e�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������A��^�U���%�6�;�!�;�l�G�������C9��Y�����6�d�h�4��4�(�������C��D��*���
�|�|�u�?�3�W���Y���F�N�����f�u�h�2�'�;�(��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���}�%�6�;�#�1����H����C9��N�����-�!�:�1��8�(��A����C9��Y�����e�u�;�u�6�����&����P9��
N��*���
�&�$���-�(���J����lR���]´�
�:�&�
�8�4�(���Y����VO��Y
�����6�;�d�'�0�o�D���Y����\��h��*���4�1�}�%�4�3��������[��G1�����0�
��%�g�.�߁�
����O�C�����u�u�u�u�w�}�W���&����[��E�� ��e�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�=�u�0�#�.����Q����`9��ZG��ʡ�0�&�4�0�:�>����Y��ƹF��G1��*���
�&�<�;�'�2�W�������@F��G1��*���y�4�
�0�w�-����	����]9��1��E���%�'�2�%�>�8�(���&������D�����c�f�u�-�#�2�ށ�����l�������6�0�
��'�m����&����OǻN�����_�u�u�u�w�<�Ͽ�&����@��Dd��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����R��^	�����b�|�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����@��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��D���8�e�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��P^�����u�k�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����C��R ��ڊ�!�|�4�1�9�)�_�������l
��h^��U���!�:�1�
�"�e�A���P�ƭ�WF��CF�����;�!�9�2�4�l�JϿ�&����C��R ��ڊ�!�|�|�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����CV��C	�����g�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��D���8�g�h�u�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����V��G�����e�<�d�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����l ��h\�����;�!�}�%�4�3��������[��G1�����<�0�
�%��)�^���P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�!�g�3�:�n�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���%�
�!�g�1�0�D��Y���F�N��U���u�%��
�$�}�JϿ�&����CV��C	�����a�_�u�u�w�}�W�������C9��h��*���f�3�8�a�j�}�W���Y���F�N�����
�&�u�h�6��#���I����9��Z1����u�u�u�u�w�5�Ͽ�&����G^��D��U��_�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F���ʺ�=�'�u�k�w�}�W���Y���F���;���&�u�h�w���/��Y���F��Y
�����_�u�u�;�w�/����B���F������u�&�<�;�'�2����Y��ƹF��G1�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�O������F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ׁ�
����O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�:�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�3�8�����Ƽ�\��D@��X���u�4�
�1�2�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����|�u�u�7�0�3�W���Y����UF�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��[��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������,�4�&�2�w�/����W���F�V�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O����ߊu�u�u�u�w�}�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�'�4�.�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Z�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lV��Y������b�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����H���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�9�>����0�ѓ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�d�u�&�>�3�������KǻN�����2�7�1�d�d�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�e� �$�<����&˹��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����f�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l3��T�����m�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����T��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����f��V��4���
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e� �&�6�8�6���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����d�4�&�2�w�/����W���F�V�����1�
�f�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�;�6�;�9�>��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�֓�]��[��<��
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������V��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�]��[��<��
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e� �&�6�8�6���H����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����a�u�&�<�9�-����
���9F������7�1�d�l�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�e� �&�6�8�6���K����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����f��V��4���g�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����S��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����f��V��4���f�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���A�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�;�4�1����H����l��G�U���0�1�%�:�2�.�}�ԜY�����D�����d�g�u�&�>�3�������KǻN�����2�7�1�d�e���������PF��G�����4�
�<�
�$�,�$���	ù��TV��D��Yʰ�<�6�;�d�1��Cف�K���F��P��U���u�u�u�u�w�}��������W9��]��H���4�
�:�&��2����Y�ƭ�l��h�����
�%�
�!�g�;���Y����]	�������!�9�d�e�j�8�����ד�F9��1��\���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�l�@���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�g���������R��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�c�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����0��
�a�6�����B����������n�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�C���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����0��
�`�6�����Y����V��=N��U���u�u�u�u�w�-��������P�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������lW��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�`�<����Y����V��C�U���4�
�<�
�3��F؁�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(߁�	����l�N�����u�u�u�u�w�}�W�������T9��S1�B��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�g�4�$�:�W�������K��N�����<�
�1�
�e�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���Y���R��d1����1�"�!�u�~�`��������_��G�U���0�1�%�:�2�.�}�ԜY�����D�����g�c�4�&�0�}����
���l�N��*���
�1�
�g��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����T��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�5�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�g�`�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b��g�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Aʴ�&�2�u�'�4�.�Y��s���R��^	�����a�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*݊�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����M���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b��d�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��]�����;�%�:�0�$�}�Z���YӇ��@��U
��G���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��7���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�E��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����P��V�����'�6�&�{�z�W�W���	����l��h\�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h,��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��k�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������`�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�g�f�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����A�ƭ�@�������{�x�_�u�w�-��������V��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ѓ�lQ��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F�� 1��B���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����g�l�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��hV�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��d�W�������A	��D�X�ߊu�u�%�&�0�?���A����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@���@����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����q9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�f�`�<����Y����V��C�U���4�
�<�
�3��G؁�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u���(�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��E���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��V��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�d�w�.����	����@�CךU���%�&�2�7�3�n�A���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�`��Fށ�	����l�N�����u�u�u�u�w�}�W�������T9��S1�C��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�N����9��h��\��u�u�0�1�'�2����s���F������7�1�f�`�6�.��������@H�d��Uʴ�
�<�
�1��o�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
���E���&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�f�u�$�4�Ϯ�����F�=N��U���&�2�7�1�d�i��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�b��l�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��]�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����;����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�f�f�4�$�:�W�������K��N�����<�
�1�
�c���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
��i������ƹF��R	�����u�u�u�u�w�}�W���
����W��]��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�&�ғ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�`�u�&�>�3�������KǻN�����2�7�1�f�e�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�b��f��������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@���Hƹ��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����f�d�4�&�0�}����
���l�N��*���
�1�
�c��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&���� P��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�:�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�e�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�l��d�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Lʴ�&�2�u�'�4�.�Y��s���R��^	�����b�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ӊ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����N���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�l��e�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��V�����;�%�:�0�$�}�Z���YӇ��@��U
��F���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��8���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�D��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&���� _��V�����'�6�&�{�z�W�W���	����l��h]�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h#��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��d�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������a�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�
9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�a�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����HӇ��Z��G�����u�x�u�u�6���������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�I����P��S/��E���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�i�W��Qۇ��P	��C1�����d�h�%�e��.����8����R��[
�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�@ʴ�&�2�u�'�4�.�Y��s���R��^	�����d�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ӊ�
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����H���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�l��a�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��Z�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��8���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�C��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����U��V�����'�6�&�{�z�W�W���	����l��hZ�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h#��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��n�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������m�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�
9��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�e�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������W��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ߓ�lW��V�����u�u�7�2�9�}�W���Y���F������7�1�a�d�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hW��*���4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���IӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ʹ��W��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�c�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��Dۊ�%�#�1�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�@����9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�a�l�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h#��G���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�b�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��z1�*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��O���
������T��[���_�u�u�%�$�:����M�ѓ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����4����R��[
��U���7�2�;�u�w�}�W���Y�����D�����a�b�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����l_��h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�i�AϿ�
����C��R��U���u�u�4�
�>�����@Ź��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ց�&�ӓ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����l�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�
9��[�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��m�����Ƽ�\��D@��X���u�4�
�<��9�(�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�m�"�������z9��V�����u�u�7�2�9�}�W���Y���F������7�1�`�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����0��
�
�'�+����s���V��G�����_�_�u�u�z�<�(���&����R��V�����'�6�&�{�z�W�W���	����l��h[�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�a�u�h��-��������lW���6���&�}�u�:�9�2�D���s���V��G�����_�_�u�u�z�<�(���&����S��V�����'�6�&�{�z�W�W���	����l��h[�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�`�u�h��-��������lW���6���&�}�u�:�9�2�C���s���V��G�����_�_�u�u�z�<�(���&����P��V�����'�6�&�{�z�W�W���	����l��h[�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�c�u�h��-��������lW���6���&�}�u�:�9�2�F���s���V��G�����_�_�u�u�z�<�(���&����_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lV��Y������g�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����L���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�e� �$�<����&����l��G�U���0�1�%�:�2�.�}�ԜY�����D�����c�f�4�&�0�}����
���l�N��*���
�1�
�b��.����	����	F��X��´�
�!�'�y�'�m�"�������z9��V�����;�&�2�u����������lW��G1�����
�<�y�%�g���������9��h��*���&�2�u�
��3��������l��A�����<�y�%�e��.����8����R��[
�����2�u�
�
�9�>����0�ӓ�C9��S1��*���y�%�e� �$�<����&Ź��l��h�����u�
�
�;�4�1����N����E
��^ �����%�e� �&�6�8�6���&����_��Y1�����
�
�;�6�;�9�>�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�e� �&�4�2��(�������W9��h��Yʥ�b��e�4��1�(���
���C9��u1�����9�
�;�&�0�}�(؁�&����l��h�����u�
�
�
��-��������TJ��hY��*ފ�%�#�1�<��4�[Ϯ�N����l��A�����<�y�%�b��k��������l��N��B���b�4�
�9��3����Y����q9��V�����;�&�2�u���(ց�	����l��D��U���
�
�e�4��1�(���
���C9��u1�*���#�1�<�
�>�q����;����R��[
�����2�u�
�
��n��������l��N��B���d�
�%�#�3�4�(���UӖ��l$��1��*���
�;�&�2�w��(���&����_��Y1�����
�
�
�
�'�+����&������h#��*���#�1�<�
�>�q����4�Փ�C9��S1��*���y�%�l��c�<�(���&����Z�G1��8���4�
�9�
�9�.����&ʹ��9��h��*���&�2�u�
���(�������]9��PB��*ӊ�
�
�%�#�3�4�(���UӖ��l+��h�����<�
�<�y�'�d�:��&����_��Y1�����
�
�
�d�6���������F��1��D؊�%�#�1�<��4�[Ϯ�@���� 9��h��*���&�2�u�
���C���&����Z��^	�����d�
�%�!�9������ƹF��R	�����u�u�u�u�w�}�W���
����W�� ]��H���%�l��e�6���������[��G1�����9�2�6�e�w�/�_���&����R��[
�����2�h�4�
�8�.�(�������	����*���
�%�#�1�>�����Y����\��h�����|�:�u�%�n��D���&����Z��^	��U���6�;�!�9�0�>�G����μ�
9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�
�'�+����&����F��h�����:�<�
�|�8�}����4�Г�C9��S1��*���u�u�%�6�9�)�������\�G1��8���4�
�9�
�9�.�������]��[����u�'�}�
���(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l+��h�����<�
�<�u�w�-��������Z��N��U¥�l��d�
�'�+����&����F��h�����:�<�
�|�8�}����4����R��[
�����2�h�4�
�8�.�(�������	����*���g�4�
�9��3����DӇ��P	��C1�����e�u�'�}���(�������W9��h��U���%�6�;�!�;�:���Y���C9��z1�*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�l��f���������@��
N��*���&�
�:�<��t����	�ѓ�lV��G1�����
�<�u�u�'�>��������lV�X������d�4�
�;���������C9��Y�����6�e�u�'���(���&����_��Y1����4�
�:�&��2����PӉ����h,��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b��c�<�(���&����Z������!�9�2�6�g�}����&Ĺ��9��h��*���&�2�h�4��2��������O��EN��*݊�
�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�j�5�������W9��h��U���%�6�;�!�;�:���Y���C9��u1�����9�
�;�&�0�`��������_	��T1�U���}�
�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�N����9��h��*���&�2�h�4��2��������O��EN��*݊�
�d�4�
�;���������C9��Y�����6�e�u�'���(���K����E
��^ �����u�%�6�;�#�1����I�ƣ�N�� 1��Dي�%�#�1�<��4�W���	����@��X	��*���:�u�%�b��l�(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l$��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�;�6�;�9�>�������W9��h��U���%�6�;�!�;�:���Y���C9��b ������
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G���
����W'��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�;�6�;�9�>�������W9��h��U���%�6�;�!�;�:���Y���C9��b ������
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G���
����W'��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�;�6�;�9�>�������W9��h��U���%�6�;�!�;�:���Y���C9��b ������
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G���
����W'��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�;�6�;�9�>�������W9��h��U���%�6�;�!�;�:���Y���C9��b ������
�e�4��1�(���
�����T�����2�6�e�u�%�u�(߁�����V��h_�����9�
�;�&�0�`��������_	��T1�U���}�
�
�;�4�1����H����l��h�����h�4�
�:�$�����&����AF��h^�����9�1��d��-��������TF�V�����
�:�<�
�~�2�WǮ�I����P��S/��Dފ�%�#�1�<��4�W���	����@��X	��*���:�u�%�e��.����8����l��A�����<�u�u�%�4�3��������F��F��*���'�u�u�%�4�3��������O��N�����%�:�0�&�]�W�W���TӇ��@��U
��C��4�&�2�u�%�>���T���F��h��*���
�b�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����C9��P1����f�_�u�u�2�4�}���Y���F�N�����<�
�1�
�`�}�J�������]��[����h�4�
�<��.����&����U��G�����:�}�%�&�0�?���J����F�R �����0�&�_�_�w�}�ZϿ�&����Q��V�����;�%�:�0�$�}�Z���YӇ��@��U
��CҊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��h^�����9�1��f�6�����Y����V��=N��U���u�u�u�u�w�-��������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�g��������� 9��h��\��u�u�0�1�'�2����s���F������7�1�b�u�$�4�Ϯ�����F�=N��U���&�2�7�1�`���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�9�>����0�ғ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����b�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l3��T�����a�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����A����@��YN�����&�u�x�u�w�<�(���&����U��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��M��i�u�4�
�8�.�(���&���R��d1����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����A�ƭ�@�������{�x�_�u�w�-��������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ù��@��R
��*ߊ�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��A��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�;�6�9�3��B���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��D���&�<�;�%�8�8����T�����D�����l�e�4�&�0�����CӖ��P�������1�
�0�
�g�e�W���
����@��d:��ڊ�!�e�3�8�f�}��������G��G����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�d�w�`�_ǻ�����WW��R	��E��h�4�
�:�$��ށ�PӇ��N��h�����:�<�
�u�w�-��������`2��G^�����3�8�d�u�9�}��������_	��T1�Hʴ�
�0�
�%�#�3�������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�@ʴ�&�2�u�'�4�.�Y��s���R��^	�����d�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�}�J���	����@��A_��U���%��
�&��}�������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�U���<�;�%�:�2�.�W��Y����C9��P1����
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���6�9�1��a�<�(���P�����^ ךU���u�u�u�u�w�}��������l_��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m�"�������z9��V�����n�u�u�0�3�-����
��ƓF�C�����2�6�0�
��-�G���ù��^9��V�����'�6�&�{�z�W�W���	����l��F1��*���
�!�e�3�:�l��������\������}�%�&�2�5�9�B��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��E���8�d�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���%�e�&�2��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ڊ�!�d�3�8�e�<����Y����V��C�U���4�
�<�
�$�,�$���	ù��TW��D��*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�m�m�u�?�3�}���Y���F�V�����&�$��
�'���������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l��1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���&����l ��h]�����;�%�:�0�$�}�Z���YӇ��@��T��*���%�e�&�2��.�(܁�
����l��TN����0�&�4�
�>�����M��ƹF��R	�����u�u�u�3��-��������V�C��U���u�u�u�u�w�<�(���&����l5��G�����
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�%�
�#�o����J���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���e�&�2�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l��1�����4�&�2�
�%�>�MϮ�������D�����`�`�_�u�w�8��ԜY���F��F��*���
�1�
�`�~�)����Y���F�N�����2�6�0�
��-�G�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������C��D��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ד�@�������%�:�0�&�w�p�W�������T9��R��!���d�3�8�e�6�.���������T��]���&�2�7�1�e�t�W�������9F�N��U���}�%�&�2�5�9�E�������9F�N��U���u�%�&�2�4�8�(���
�ד�@��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��M���8�`�4�&�0�����CӖ��P�������7�1�l�`�]�}�W������F�N��U´�
�<�
�1��l�^Ϫ���ƹF�N��U���%�&�2�6�2��#���A����lS�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����G^��D��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��O�����
� �m�c�'�}�J���[ӑ��]F��{1��*���
�:�%�`�'�4����K����[��G1�����9�`�d�|�2�.�W��B��� ��[�����:�%�d�
��5�(���H����CU�
NךU���u�u�
�
������ӑ��]F��R�����3�
�l�
�e�m�W���H����_��=N��U���u�0�
�8�f����L����l�N��*����'��:��i�F�������T��h�I���u�u�u�u�'�d�:�������TF��R �����!�%�l�3��l�C���Q���A��N�����u�u�u�u�$�1����L����T��h����u�u�u��9�9�(����Փ�F9��^��D��u�!�
�:�>�����۔��Z��D������-� �,�"��(���&����J��G����u�u�u��9�9�(�������@9��h_�A���u�h�&�1�;�:��������A��M�����1�<�
������&¹��T9��]��F���n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������l^��h�����2�
�'�6�m�-����
ۇ��A��G�����%�
�!�y�6�����
����g9��1��ي�&�
�y�4��4�(�������C��D��*���
�y�4�
�2���������l��N��*����'��:��i�G�������lT��B��&���
�:�
�:�'�l�(ށ�����T9�� V��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��4�(�������C��D��*���
�|�4�1��-��������Z��S�����2�%�<�0��-�(���P����[��=N��U���u�u�u�'��(�O���	��� ��[�����:�%�d�
��5�(���&����l�N��Uʰ�&�3�}�}�'�>��������lW������%�<�0�
�'��������R��X ��*���<�
�u�u�'�.��������l��h��F���8�a�|�u�?�3�}���Y���F�P�����f�
�e�i�w���������\��1�����'�2�g�e�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�e�G���Y���k>��o6��-���������/���!����l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����3�
�f�
�f�a�W���&����9l�N�U���
� �m�a�4�}����Ӗ��P��N����u�'�
� �o�i����
����l��TN����0�&�4�
�2�}��������B9��h��*���g�3�8�f�w�%����¹��T9��V����<�
�&�$���߁��Փ�@��N��*���
�&�$���-�(���H����lT�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W�������\��h��*��m�h�4�
�8�.�(���&����]�V�����
�:�<�
�w�}��������B9��h��*���d�3�8�g�~�2�W���	����@��X	��*���u�%�&�2�4�8�(���	�֓�G��Q��F���;�u�}�-�#�2�ށ����� ^������!�9�d�e�~�}��������\��h��*��m�h�4�
�8�.�(���&����]�V�����
�:�<�
�w�}��������B9��h��*���f�3�8�a�~�t�W������F�N��Uʲ�%�3�
�f��8�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F�	��*���m�a�6�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�'��(�O���	�ƭ�@�������{�x�_�u�w�/�(���A�ғ�9��D��*���6�o�%�:�2�.��������V��c1��E���2�
�&�
�{�<�(���&����V��G^�����3�
�:�0�#�/�(܁�����9��N��*���
�&�$���-�(���H����lT�Q=�����!�'�
�a�$�;�(��M����9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�0�
�%�#�3���������Yd��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	����
����U��G�����u�u�u�u�w�}�W���YӁ��l ��]�����h�3�
�:�2�)����M����F9��Z��D�ߊu�u�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����CV��C	�����g�|�!�0�w�}�W���Y���F�	��*���m�a�%�u�j�;�(�������^9��Q��F���%�n�u�u�w�}�W�������9F�N��U���u�u�u�'��(�O���	���D��o6��-���������/���!����kD��N��U���u�u�0�1�>�f�W���Y����_��=N��U���u�u�u�'��(�O���	���D��o6��-���������/���!����kD��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʼ�
�<��'��2�(ځ�&����G9��h_�G���u�h�}�8��(�O���	�ƣ���T�����a�d�n�u�w�4�(���?����\	��1��D���
�g�a�%�w�`��������l��C�� ���2�0�}��;���������l��h��M���%�|�~� �$�:����	����@��A[��\��_�u�u�x�>���������C9��G�����g�
�a�4�$�:�W�������K��N�����<��'��8��(���&����T��1�����
�'�6�o�'�2��������l ��h"�����'�2�m�m�w�%����¹��T9��V����<�
�&�$���߁��֓�@��N��*���
�%�!�;�'�m���Y����Z9��E1�����
�
�
�0��l�O�ԜY�Ʈ�T��N��U���<�u�}�0�>�>��������U��
N��*���&�
�#�
�~�<����	����@��X	��*���u�%�&�2�4�8�(���	�֓�G��Q��D���;�u�4�
�8�.�(�������F��h��*���!�;�%�e�>�l�^������F�N��U���<�
�<��%�����&����U��\��A��u��9�
�8�����L�ד�l��h\�M�ߊu�u�u�u�;�8�}���Y���F�^"�����'��:�
��5�(���A�ԓ�F������:�
�:�%�b�/���A���F�N��ʼ�n�_�u�u�9�}����
��ƓF�^9��&����!�d�
��(�F��&���F��S1�����#�6�:�}�9�4��������_T��Q��D���%�|�x� �$�:��������Q��B1�F؊�f�|�_�u�w�
���� ����@9��h_�C���u�h�&�1�;�:��������F��P ��]����9�
� �n�o����Tӓ��Z��SF�����d�
� �d�f��D���s���]��R�*���l�m�%�u�j�W�W���Y�Ƽ�9��1��*���u�=�;�}�2���������l��G��U��|�0�&�u�w�}�W���	�ѓ�lW��^ ����u�u�;�"�2�l�(���@�ғ� F�d��U���u�;�"�0�`�;�(��&����[�������
� �l�a�'�u�^��^���V
��d��U���u�;�"�0�o�;�(��&����F�Y����
� �d�e��n�K���Y���F��R��ӊ� �l�g�%�w�5��������WT��B1�M���}�|�h�r�p�}����s���F�Y����
� �l�m�'�f�W�������_W��Q��E���%�u�h�_�w�}�W�������W��B1�A���u�=�;�}�%�>��������9��^��H��r�u�9�0�]�}�W���Y����V
��h��D��
�f�_�u�w�8�$���M����W��h�I���u�u�u�u�'�m�"�������z9��^ �����=�;�}�0��0�Fց�����9��^��H��r�u�9�0�]�}�W���Y����f��V��4���f�<�
�<�l�}�Wϰ�����9��h_�G���u�h�_�u�w�}�W���&����R
��v'��D���
�<�u�=�9�u��������U��^�����|�h�r�r�w�1��ԜY���F��1�����0��
�
�9�.��ԜY�Ƣ�D5��X�� ��a�
�f�i�w�}�W���YӖ��l3��T�����b�<�
�<�w�5��������CW��Q��E���%�}�|�h�p�z�W������F�N��E���&�4�0����������F��@=��D݊� �d�`�
�d�a�W���Y�����h;�����1��f�<��4�W����ο�_9��G_�����e�m�%�}�~�`�P���Y����l�N��Uʥ�e� �&�4�2��(�������T]ǻN�����9�m�3�
�f�o����D���F�N�����d�
� �d�e��Dϩ�����A9��Y
�����d�c�%�}�~�`�P���Y����l�N��Uʻ�"�0�d�
�"�l�D݁�J���F��@=��Dӊ� �d�b�
�d�a�W���Y�����d��C���
�d�a�%�w�5��������WR��B1�@ڊ�g�e�u�u�f�t����Y���F� ��&���b�3�
�d�a�-�L���Yӈ��`��h��L���%�u�h�_�w�}�W���&ù��@��R
��*���<�
�<�u�?�3�_���&����l ��V�����|�h�r�r�w�1��ԜY���F��1�����0��
�
�9�.��ԜY�Ƣ�D5��^�� ��m�
�f�i�w�}�W���Yӈ��`��1��*��g�%�u�=�9�u�����ӓ�F9�� ^��G��u�u�d�|�2�.�W���Y�����d��L���
�d�c�%�l�}�Wϰ�����9��h_�G���u�h�_�u�w�}�W���&����Z��^	�����}�0�
�8�f����Hǹ��V�
N��R���9�0�_�u�w�}�W���&����l��D�����u�0��9�e�;�(��A����[�N��U���%�b��d��3����������h��D݊� �d�e�
�e�m�W���H����_��=N��U���u�
�
�
��3����s���]��R�*���d�e�
�f�k�}�W���Y����lQ��hY�����2�"�0�u�$�1����L����V��h�E���u�d�|�0�$�}�W���Y����lQ��h[�����2�_�u�u�2���������V��N�U���u�u�u�%�`��D���&����D��F�����%�f�3�
�g�e����P���A�R��U���u�u�u�%�`��Fځ�����l�N�����g�
� �d�f��D��Y���F� ��&���d�3�
�d�e�-�W����Σ�l��SV�� ��g�
�g�e�w�}�F�������9F�N��U����9�g�3��l�O���B�����d��C���
�g�a�%�w�`�}���Y���]��R�*���d�e�
�f� �8�WǱ�&����9��h_�E���}�|�h�r�p�}����s���F�Y����
� �d�d��n�}���Y����V
��h��D��
�f�i�u�w�}�W�������_T��Q��G���%�u�=�;��/����L����W��h�E���u�d�|�0�$�}�W���Y����V��[\�����g�a�%�n�w�}�����ԓ�F9��1��U��_�u�u�u�w��(�������r/��h�����"�0�u�&�;�)�ہ�����l��G��U��|�0�&�u�w�}�W���	�֓�]��[��<���<�
�<�n�w�}�����Փ�F9��1��U��_�u�u�u�w��(�������r/��h�����"�0�u�&�;�)����&����CT�N��R��u�9�0�_�w�}�W���&ù��@��R
��*���<�
�<�n�w�}�����ғ�F9��1��U��_�u�u�u�w�8�$�������9�������'�6�;�
�"�d�C���Q���A��N�����u�u�u�u�9�*��������9��d��Uʻ�"�0�`�3��h�(��E��ƹF�N�����9�
� �l�e�-�W����Σ�l��S\�� ��m�%�}�|�j�z�P������F�N�����0�f�3�
�d��D�ԜY�Ƣ�D5��1��*��
�f�i�u�w�}�W�������_R��B1�E���u�=�;�}�%�>��������9��^��H��r�u�9�0�]�}�W���Y����V
��Q��@ފ�f�_�u�u�2��؁�����l��S��U���u�u�%�b��m�����ƻ�V�D�����
� �m�g�'�u�^��^���V
��d��U���u�%�b��f��������F��@=��M���
�b�
�f�k�}�W���Y����lQ��h_�����<�u�=�;��8�(���A����^��G\��\��r�r�u�9�2�W�W���Y�Ƽ�9��1��*���n�u�u�;� �8�N���&����CU�
NךU���u�u�
�
������ӑ��]F��R�����3�
�c�
�e�m�W���H����_��=N��U���u�
�
�
��3����s���]��R�� ��m�%�u�h�]�}�W���Y����f��V��4���
�;�&�2� �8�Wǭ����� 9��hV�*��e�u�u�d�~�8����Y���F��h^�����9�1��d��3����s���\��X ��*���l�c�%�u�j�u�����ޓ�F9��1��U���&�9�!�%��(�O���	����F�X�����
� �l�m�'�}�J�������CR��B1�M���u�'�&�9�#�-�(���A�ԓ�O��N�����:�1�
� �n�e����D�Σ�l��S1��*��
�g�:�u�%�>��������9��UךU���'�6�;�a�1��F���	���N��[1�����3�
�e�e�'�}�ϭ�����R��B1�Mފ�g�n�u�u�8�����&����Q��G\��H���'�6�;�m�1��F���	�ƣ�	��T��L���
�d�m�%�~�W�W�������W^��B1�G܊�g�i�u�&�;�)��������R��N��U���
�8�d�
�"�l�Gׁ�K��ƹF��E1�����3�
�d�m�'�}�J�������CW��Q��D���%�u�'�&�;�)��������
P��G�U���:�
�:�1�1��Gہ�K�����h��F���
�l�
�g�8�}�����ד�F9��1��\�ߠu�u�x�u����������lV��G1�����
�<�u�&�>�3�������KǻN��*ڊ�;�6�9�1��m��������l��h�����%�:�u�u�%�>����&ù��@��R
��*ڊ�%�#�1�u����������lV��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��v'��*���#�1�|�!�2�}�W���Y���F��h^�����9�1��e�6���������Z�G1�� ���4�0��
��-����s���F�R��U���u�u�u�u�w�-�G���
����W'��1��*���
�;�&�2�k�}�(߁�����V��h^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l3��T�����e�<�
�<�w�.����	����@�CךU���
�
�;�6�;�9�>�������T9��D��*���6�o�%�:�2�.����,����_��~1�U���
�;�6�9�3��G�������lV��Y������e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��b ������
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�;�6�;�9�>�������TF���*���6�9�1��g�W�W���Y�Ʃ�@�N��U���u�u�%�e��.����8����Z��^	��Hʥ�e� �&�4�2��(߁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(�������W9��h��U���<�;�%�:�2�.�W��Y����lV��Y������d�
�%�!�9��������@��h����%�:�0�&�'�m�"�������z9��h�����u�
�
�;�4�1����Hù��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�m�"�������z9��h�����|�!�0�u�w�}�W���Y����lV��Y������d�
�%�!�9���������h;�����1��d�
�'�+��ԜY���F��D��U���u�u�u�u�'�m�"�������z9��h�����<�
�<�u�j�-�G���
����W'��^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l3��T�����d�
�;�&�0�<����Y����V��C�U���%�e� �&�6�8�6���I����@��V�����'�6�o�%�8�8�Ǯ�I����P��S/��D���%�e� �&�6�8�6���I����TJ��h^�����9�1��d��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���6�9�1��f���������[��=N��U���u�u�u�
��3��������9��h��U��%�e� �&�6�8�6���I���F�N�����u�u�u�u�w�}����,����_��~1�*���&�2�i�u����������lW��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�"�������z9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��Fށ�	����l��D�����2�
�'�6�m�-����
ۖ��l3��T�����d�
�%�#�3�}�(߁�����V��h_�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l3��T�����d�
�%�#�3�t����Y���F�N��U���
�;�6�9�3��Fށ�	����l��D��I���
�
�;�6�;�9�>��&����_��N��U���0�&�u�u�w�}�W���YӖ��l3��T�����d�
�%�#�3�4�(���Y����lV��Y������d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��l�(���
����@��YN�����&�u�x�u�w�-�G���
����W'��_�����2�4�&�2��/���	����@��h^�����9�1��d�{�-�G���
����W'��_�����u�
�
�;�4�1����H¹��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�9�>����0����R��[
��U���;�_�u�u�w�}�W���&ù��@��R
��*���<�
�<�u�j�-�G���
����W'��_�U���u�u�0�&�w�}�W���Y�����h;�����1��d�
�9�.���Y����f��V��4���d�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l3��T�����d�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������lW��V�����;�&�2�4�$�:�(�������A	��D��*ڊ�;�6�9�1��l�(������C9��b ������
�g�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ڊ�;�6�9�1��l�(��������YNךU���u�u�u�u����������lW��V�����;�&�2�i�w��(�������r/��1��*���n�u�u�u�w�8����Y���F�N��*ڊ�;�6�9�1��l�(�������]9��PN�U���
�;�6�9�3��F݁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��3��������9��h��U���<�;�%�:�2�.�W��Y����lV��Y������d�
�;�$�:��������\������}�
�
�;�4�1����H����lV��Y������d�
�'�0�}�(߁�����V��h_�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��v'��G���
�9�|�u�?�3�}���Y���F�G1�� ���4�0��
�e�4�(���Y����lV��Y������d�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�;�6�;�9�>��&����Z�
N��E���&�4�0���o����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��l�(�������]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���f�4�
�9��3��������]9��X��U���6�&�}�
��3�������� 9��h��Yʥ�e� �&�4�2��(�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��3�������� 9��h��\���=�;�_�u�w�}�W���Y����f��V��4���f�4�
�9��3����E�Ƽ�9��D�����
�f�4�
�;�f�W���Y����_��=N��U���u�u�u�
��3�������� 9��h��*���&�2�i�u����������lW��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��F܁�����l��^	�����u�u�'�6�$�u�(߁�����V��h_�U���
�;�6�9�3��F܁����C9��b ������
�f�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����0��
�f�6�����Y����l�N��U���u�%�e� �$�<����&�Փ�]9��PN�U���
�;�6�9�3��F��Y���F��[�����u�u�u�u�w��(�������r/��1��*���u�h�%�e��.����8����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��3��������9��h��*���&�2�4�&�0�}����
���l�N��E���&�4�0���i��������l��h�����%�:�u�u�%�>����&ù��@��R
��*���4�
�9�y�'�m�"�������z9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��@��R
��*���4�
�9�|�w�5��ԜY���F�N��E���&�4�0���i��������l��R����� �&�4�0���C���&����9F�N��U���0�_�u�u�w�}�W���&ù��@��R
��*���4�
�9�
�9�.���Y����f��V��4���a�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
�c�4�(���Y����T��E�����x�_�u�u����������lW��^ �����&�<�;�%�8�}�W�������C9��b ������
�a�u����������lW��G��Yʥ�e� �&�4�2��(�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e� �&�6�8�6���M����E
��N�����u�u�u�u�w�}����,����_��~1�*���&�2�i�u����������lW��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��D�����
�a�<�
�>�}�JϮ�I����P��S/��Dފ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e��.����8����l��A�����<�
�&�<�9�-����Y����V��G1�� ���4�0��
�b�<�(���UӖ��l3��T�����d�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�� ���4�0��
�b�<�(���P�Ƹ�V�N��U���u�u�%�e��.����8����l��A�����<�u�h�%�g���������S��G1���ߊu�u�u�u�;�8�}���Y���F�G1�� ���4�0��
�b�<�(���&����Z�
N��E���&�4�0���h��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�e� �$�<����&�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���`�<�
�<��.����	����	F��X��¥�e� �&�4�2��(��Y����f��V��4���`�%�0�y�'�m�"�������z9��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G���
����W'��[�����1�|�!�0�w�}�W���Y�����h;�����1��d�
�9�.���Y����f��V��4���`�_�u�u�w�}����s���F�N����� �&�4�0���B���&����[��h^�����9�1��d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
��-��������TF��D��U���6�&�{�x�]�}�W���&����R
��v'��*���#�1�<�
�>���������PF��G�����%�e� �&�6�8�6���&����_�G1�� ���4�0��
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e� �&�4�2��(ށ�	����O��_�����u�u�u�u�w��(�������r/��h�����<�
�<�u�j�-�G���
����W'��1��*���n�u�u�u�w�8����Y���F�N��*ڊ�;�6�9�1��l��������l��R����� �&�4�0���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�9�>����0�ד�]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���
�;�&�2�6�.���������T��]���
�;�6�9�3��F���&ù��@��R
��*ۊ�'�2�u�
��3��������l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g���������9��h��\���=�;�_�u�w�}�W���Y����f��V��4���
�;�&�2�k�}�(߁�����V��h_�U���u�u�0�&�w�}�W���Y�����h;�����1��d�<��4�W��	�֓�]��[��<���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�֓�]��[��<���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e��.����8����R��[
�����2�4�&�2��/���	����@��h^�����9�1��g�6����	�֓�]��[��<���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h;�����1��g�4��1�^������F�N��U���%�e� �&�6�8�6���&����_��Y1����u�
�
�;�4�1����K����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��D�����
�
�%�#�3�4�(���Y����lV��Y������g�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��E���&�4�0�������Ӈ��Z��G�����u�x�u�u�'�m�"�������z9��^ �����&�<�;�%�8�}�W�������C9��b ������
�y�%�g���������9��R	���� �&�4�0���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�;�6�9�3��E���&����F��R ��U���u�u�u�u�'�m�"�������z9��^ �����h�%�e� �$�<����&��ƹF�N�����_�u�u�u�w�}�W���&����R
��v'��*���&�2�i�u����������lT��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u����������lU��G1�����
�<�u�&�>�3�������KǻN��*ڊ�;�6�9�1��n��������l��h�����%�:�u�u�%�>����&ù��@��R
��*ي�%�#�1�u����������lU��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��v'��*���#�1�|�!�2�}�W���Y���F��h^�����9�1��f�6���������Z�G1�� ���4�0��
��-����s���F�R��U���u�u�u�u�w�-�G���
����W'��1��*���
�;�&�2�k�}�(߁�����V��h]�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l3��T�����f�<�
�<�w�.����	����@�CךU���
�
�;�6�;�9�>�������T9��D��*���6�o�%�:�2�.����,����_��~1�U���
�;�6�9�3��D�������lV��Y������f�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��b ������
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�;�6�;�9�>�������TF���*���6�9�1��d�W�W���Y�Ʃ�@�N��U���u�u�%�e��.����8����Z��^	��Hʥ�e� �&�4�2��(܁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(ہ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�g���������9��h��Yʥ�e� �&�4�2��(ہ�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�e��.����8����R��[
��U���;�_�u�u�w�}�W���&ù��@��R
��*ފ�%�#�1�<��4�W��	�֓�]��[��<���4�
�9�n�w�}�W�������9F�N��U���u�
�
�;�4�1����M����E
��^ �����h�%�e� �$�<����&ǹ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������r/��h�����4�&�2�u�%�>���T���F��1�����0��
�
�9�.����
����C��T�����&�}�
�
�9�>����0���C9��b ������
�
�'�0�}�(߁�����V��hZ�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����,����_��~1�����9�|�u�=�9�W�W���Y���F��1�����0��
�
�9�.���Y����f��V��4���n�u�u�u�w�8����Y���F�N��*ڊ�;�6�9�1��i���������h;�����1��a�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h;�����1��`�4��1�(���
����@��YN�����&�u�x�u�w�-�G���
����W'��1��*���
�;�&�2�6�.���������T��]���
�;�6�9�3��B���&������h;�����1��`�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ڊ�;�6�9�1��h�������G��d��U���u�u�u�%�g���������9��h��*���&�2�i�u����������lS��G1���ߊu�u�u�u�;�8�}���Y���F�G1�� ���4�0��
��-��������TF���*���6�9�1��b�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�e� �&�6�8�6���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I����P��S/��@���
�<�
�&�>�3����Y�Ƽ�\��DF��E���&�4�0���q����,����_��~1�����y�%�e� �$�<����&ƹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�9�>����0�ӓ�C9��SG�����u�u�u�u�w�}�WϮ�I����P��S/��@���
�<�u�h�'�m�"�������z9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��D�����
�
�;�&�0�a�W���&����R
��v'��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��v'��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�;�4�1����O����E
��^ �����&�<�;�%�8�}�W�������C9��b ������
�
�%�!�9�W���&����R
��v'��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��D�����
�
�%�#�3�t����Y���F�N��U���
�;�6�9�3��A���&����Z��^	��Hʥ�e� �&�4�2��(ف�	����l�N��Uʰ�&�u�u�u�w�}�W���	�֓�]��[��<���4�
�9�
�9�.���Y����f��V��4���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h^�����9�1��c�>�����
������T��[���_�u�u�
��3��������l��D�����2�
�'�6�m�-����
ۖ��l3��T�����c�u�
�
�9�>����0�Г�A����*���6�9�1��a�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��E���&�4�0�����������[��=N��U���u�u�u�
��3��������l��D��I���
�
�;�6�;�9�>��s���F�R��U���u�u�u�u�w�-�G���
����W'��1��*���u�h�%�e��.����8����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e��.����8����R��[
�����2�4�&�2�w�/����W���F�G1�� ���4�0��
��-��������T9��D��*���6�o�%�:�2�.����,����_��~1�����9�y�%�e��.����8����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G���
����W'�� 1��*���|�u�=�;�]�}�W���Y���C9��b ������
�
�%�!�9���������h;�����1��b�4��1�L���Y�����RNךU���u�u�u�u����������lQ��G1�����
�<�u�h�'�m�"�������z9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*݊�;�&�2�4�$�:�W�������K��N����� �&�4�0���(���
����@��Y1�����u�'�6�&���(�������r/��N��E���&�4�0�������Y����f��V��4���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l3��T�����b�4�
�9�~�}����s���F�N����� �&�4�0���(���
���F��1�����0��
�n�w�}�W�������9F�N��U���u�
�
�;�4�1����N����@��S��*ڊ�;�6�9�1��j����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��e��������l�������%�:�0�&�w�p�W���	�֓�]��[��<���4�
�9�
�9�.����
����C��T�����&�}�
�
�9�>����0�ޓ�C9��SB��*ڊ�;�6�9�1��e��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�;�4�1����A����E
��N�����u�u�u�u�w�}����,����_��~1�����9�
�;�&�0�a�W���&����R
��v'��*���#�1�_�u�w�}�W������F�N��Uʥ�e� �&�4�2��(ׁ�	����l��D��I���
�
�;�6�;�9�>�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g���������9��h��U���<�;�%�:�2�.�W��Y����lV��Y������m�<�
�>���������PF��G�����%�e� �&�6�8�6���UӖ��l3��T�����m�%�0�y�'�m�"�������z9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(�������r/��h�����|�!�0�u�w�}�W���Y����lV��Y������m�<�
�>�}�JϮ�I����P��S/��M�ߊu�u�u�u�;�8�}���Y���F�G1�� ���4�0��
��3����E�Ƽ�9��D�����
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��D�����
�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������l_��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��E���&�4�0��������Ƽ�9��D�����
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�� ���4�0��
��-����PӒ��]FǻN��U���u�u�
�
�9�>����0�ߓ�C9��S1��*���u�h�%�e��.����8����R��[
�U���u�u�0�&�w�}�W���Y�����h;�����1��l�4��1�(���
���F��1�����0��
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�;�6�9�3��N���&����R��P �����&�{�x�_�w�}�(߁�����V��hW�����2�4�&�2��/���	����@��h^�����9�1��l�w��(�������r/��h�����
�
�;�6�;�9�>�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e� �&�6�8�6���&����_����ߊu�u�u�u�w�}�(߁�����V��hW�����2�i�u�
��3��������l�N��Uʰ�&�u�u�u�w�}�W���	�֓�]��[��<���<�
�<�u�j�-�G���
����W'��1����u�u�u�u�2�9���s���V��G�����_�u�u�%�c�����8����[��hZ�����1��7�3�2��C�������lǻN��Xʥ�a��4�0���(�������@��YN�����&�u�x�u�w�-�C�������z9��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�O������F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ׁ�
����O��_�����u�u�u�u�w��(�������lV��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����*����W'��1��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*ފ�6�9�1��f�a�W���&����V��h�����d�
�0�
�e�f�W���	�ғ�P��S/��D���h�%�a��6�8�6�������lW��Z�����a�n�_�u�w�p����*����W'��^�����1�4�&�2�w�/����W���F�G1��&���0��
�e�6�����
����l��TN����0�&�4�
�2�}��������B9��h��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��M���8�`�|�u�?�3�}���Y���F�G1��&���0��
�e�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N������4�0���m���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W���&����V��h_�I���
�
�6�9�3���������lW��E��B��_�u�u�x�w��(�������lW��V�����&�<�;�%�8�8����T�����h=������d�
�%�!�9��������\������}�%�6�y�6�����
����g9��1�����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��CV�����|�|�!�0�w�}�W���Y�����h=������d�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���*���9�1��d��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�C�������z9��R������4�0���(����H����A�� X����u�x�u�
��>����0����R��[
�����;�%�:�0�$�}�Z���YӖ��l5��[��<��
�%�#�1�6�.���������T��]���6�y�4�
�>�����*����9��Z1����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����G^��D��\���!�0�u�u�w�}�W���YӖ��l5��[��<��
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h=������d�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�%�c�����8����Z�G1��&���0��
� �1�/�F܁�&����Q��=d��U���u�
�
�6�;�9�>��&����_��D��ʥ�:�0�&�u�z�}�WϮ�M����_��~1�*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$���˹��^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����u�u�u�u�w�}�WϮ�M����_��~1�*���#�1�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӖ��l5��[��<��
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�a��6�8�6���M���C9��d�����
� �3�'�f��(���&����9l�N�U���
�6�9�1��l�(�������@��YN�����&�u�x�u�w�-�C�������z9��h�����4�&�2�
�%�>�MϮ�������T����<�
�&�$���ׁ�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C��U���u�u�u�u�w�-�C�������z9��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�M����_��~1�*���#�1�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʥ�a��4�0���B��Y����`��R
��*���3�'�d�
��8�(��B���F���*���9�1��d��-��������]F��X�����x�u�u�%�c�����8����l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�e����L���G��d��U���u�u�u�%�c�����8����l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�C�������z9��h�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�a��4�0���(�������@��YN�����&�u�x�u�w�-�C�������z9��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�O������F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ׁ�
����O��_�����u�u�u�u�w��(�������lW��G1����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����*����W'��1��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*ފ�6�9�1��e�a�W���&����V��h�����d�
�
�0��n�L�ԜY�����h=������g�4�
�;�}����Ӗ��P��N����u�
�
�6�;�9�>�������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�m�3�:�h�^������F�N��U���%�a��4�2��(݁�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�4�1����K����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�9��V��4���u�h�%�a��<����&����V��1�����c�l�_�u�w�p�W���&����V��h]�����1�4�&�2�w�/����W���F�G1��&���0��
�
�'�+����
����C��T�����&�}�%�6�{�<�(���&����l5��D�����`�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�}�W���Y���F��hZ�����1��f�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��A���4�0��
��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�C�������z9��S��*ފ�6�9�1��5�;����M�ӓ�V��\����u�x�%�a��<����&ǹ��l�������%�:�0�&�w�p�W���	�ғ�P��S/��A���
�9�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
�ޓ�@��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�_�u�u�w�}�W���&ǹ��R
��v'��*���#�1�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӖ��l5��[��<���4�
�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�
�
�6�;�9�>��E�Ƽ�9��V��4��� �3�'�d������N��ƓF�C��*ފ�6�9�1��b�<�(���Y����T��E�����x�_�u�u����������l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�e����L���G��d��U���u�u�u�%�c�����8����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w��(�������lS��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1��&���0��
�u�j�-�C�������z9��Q��*���l�'�2�c�o�W�W���T�Ƽ�9��V��4���
�%�#�1�6�.��������@H�d��Uʥ�a��4�0���(�������@��Y1�����u�'�6�&��-�������T9��R��!���m�3�8�`�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�t����Y���F�N��U���
�6�9�1��k���������T�����2�6�d�_�w�}�W������F�N��U���%�a��4�2��(ف�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W���	�ғ�P��S/��B��u�
�
�6�;�9�>�������S��h��*��n�_�u�u�z�-�C�������z9��V�����&�<�;�%�8�8����T�����h=������b�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1�����|�u�=�;�]�}�W���Y���C9��d�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��hZ�����1��b�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u����������Z�G1��&���0��
� �1�/�Fہ�O����lQ��dךU���x�%�a��6�8�6���&����_��D��ʥ�:�0�&�u�z�}�WϮ�M����_��~1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���A����lS�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9��G�����_�u�u�u�w�}�W���&����V��hV�����1�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W���	�ғ�P��S/��M���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�6�9�3��N��Y����`��R
��*���3�'�d�
�a�/���N��ƹF�N��A���4�0��
��-��������]F��X�����x�u�u�%�c�����8����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�o�;���s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P����[��=N��U���u�u�u�
��>����0�ߓ�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�i�$�������
9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��hZ�����1��7�3�2��C��&���� S��G]��H�ߊu�u�u�u�%����I����D��F�����%�
�0�
�g�n�G���Y�����RNךU���u�u�
�
�4�1��������A9��hW�����m�n�u�u�'�i�$�������Q��R��A��
� �d�`��n�K���Y���F��hZ�����1��7�3�2��C�������^��_��]���
�8�g�'�0�o�B���P���A�R��U���u�u�u�%�c�����8����U ��h_��Dڊ� �d�`�
�d�W�W���&ǹ��R
��v'�� ���'�d�
�g�1��D���	���l�N��Uʥ�a��4�0����������
9��P1�Mʢ�0�u�&�9�#�-����K����O�I�\ʰ�&�u�u�u�w�}����*����W'��U�����a�d�
� �f�h�(��s���C9��d�����
� �3�'�f��D���&����l��S��U���u�u�%�a��<����&����V��1�����c�m�"�0�w�.����	����T9��]��\��r�r�u�9�2�W�W���Y�Ƽ�9��V��4��� �3�'�d��o����J�ғ� ]ǻN��*ފ�6�9�1��5�;����M����U��Y�����h�_�u�u�w�}����M�ƻ�V�D�����
�0�
�e�e�m�W���H����_��=N��U���u�
�
�6�;�9�>�������R��1����a�_�u�u����������F ��E1�*���3�
�f�`�'�}�J�ԜY���F��1������
� �3�%�l�(�������R��_��]���
�8�a�'�0�o�A���P���A�R��U���u�u�u�%�c�����8����U ��h_��D݊� �d�b�
�d�W�W���&ǹ��R
��v'�� ���'�d�
�l�1��D���	���l�N��Uʥ�a��4�0����������P��R	��D���=�;�}�0��0�E������� N��S��D���0�&�u�u�w�}�WϮ�M����_��~1�����
�a�d�
�"�l�Oځ�J���F��1������
� �3�%�l�(ށ�����9��R�����u�u�u�'��(�O���	�ƻ�V�D�����
�0�
�e�d�m�W���H����_��=N��U���u�
�
�6�;�9�>�������R��R	��D��u�u�%�a��<����&����V��1�*���d�l�
�f�k�}�W���Y����lR��T�����7�3�0�
�c�l�(���&����D��F�����%�'�2�g�c�u�^��^���V
��d��U���u�%�a��6�8�6�������lW��W�� ��l�
�f�_�w�}�(ہ�����r/��B����
�d�3�
�c�k����D���F�N��A���4�0��
�"�;���&�Г�V��Z�����}�0�
�8�d�/���@����[�I�����u�u�u�u�w�-�C�������z9��Q��*���g�
� �d�n��D�ԜY�Ƽ�9��V��4��� �3�'�d��o����M�Փ� F�d��U���u�'�2�m�e�*����
����^��E��G��}�|�h�r�p�}����s���F�G1��&���0��
� �1�/�Fہ�M����lQ��d��Uʥ�a��4�0����������U��B1�Gڊ�f�i�u�u�w�}�WϮ�M����_��~1�����
�a�d�
�2��C������@��C��*���
�e�g�e�w�}�F�������9F�N��U���
�6�9�1��?����&�ғ�9��h_�F���n�u�u�%�c�����8����U ��h_��Gފ� �d�g�
�d�a�W���Y�����h=������7�3�0��i�Fہ�����F��R �����!�%�
�0��m�D��Y���O��[�����u�u�u�
��>����0����U��Z��F���
�a�e�%�l�}�WϮ�M����_��~1�����
�a�g�
�"�l�Dہ�J���9F�N��U���
�6�9�1��?����&�ғ�9��P1�Eʢ�0�u�&�9�#�-�(���&����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�a�3��i�@���B�����h=������7�3�0��i�Eف�����9��R�����u�u�u�
��>����0����U��Z��A���2�b�e�"�2�}��������V��Z�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�c�o�(���H����CU��N������4�0���(����Hǹ��l ��Z�*��i�u�u�u�w�}����*����W'��U�����a�d�
�0��i�W����ο�_9��G]�����e�f�e�u�w�l�^ϻ�
��ƹF�N��*ފ�6�9�1��5�;����M����U��Z����u�u�%�a��<����&����V��1�*���d�`�
�f�k�}�W���Y����V��\�����}�0�
�8�f�/���A����[�I�����u�u�u�u�w�-�C�������z9��Q��*���&�'�2�b�a�W�W���&ǹ��R
��v'�� ���'�d�
�l�1��C���	���l�N��Uʥ�a��4�0����������@9��P1�Cʢ�0�u�&�9�#�-�(���&����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�m�3��i�B���B�����h=������7�3�0��i�D߁�����
9��R�����u�u�u�
��>����0����U��\��*���
�c�u�=�9�u�����Г�V��Y�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�c�o�(���H����CU��N������4�0���(����Hǹ��l ��Z�*��i�u�u�u�w�}����*����W'��U�����g�&�'�2�`�k� ���Yە��l��1����c�}�|�h�p�z�W������F�N��A���4�0��
�"�;���&�֓�F9��W��F�ߊu�u�
�
�4�1��������A9��h]�����a�f�%�u�j�W�W���Y�Ƽ�9��V��4��� �3�'�d������O�ƻ�V�D�����
�0�
�e�d�m�W���H����_��=N��U���u�
�
�6�;�9�>�������R��1��*��c�%�n�u�w�-�C�������z9��Q��*���f�
� �d�n��D��Y���F���*���9�1��7�1�8�(���
����lQ�������0�
�8�
�2��G��I���W����ߊu�u�u�u����������F ��E1�*���3�
�a�f�'�f�W���	�ғ�P��S/�����0�
�a�f��(�F��&���FǻN��U���
�
�6�9�3���������l��R	��C���=�;�}�0��0�D������� N��S��D���0�&�u�u�w�}�WϮ�M����_��~1�����
�a�f�
�"�l�N߁�J���F��1������
� �3�%�l�(�������R��N�U���u�u�u�%�c�����8����U ��h_�����2�b�g�"�2�}��������A��^�]���h�r�r�u�;�8�}���Y���A��Z����u�
�
�6�;�9�>�������R��1��*���d�%�u�h�]�}�W���Y����`��R
��*���3�'�d�
��8�(��Y����N��[1��Ҋ�0�
�e�e�g�}�W��PӃ��VFǻN��U���
�
�6�9�3���������lU��Q��@���%�n�u�u�'�i�$�������Q��R��A��
� �d�d��n�K���Y���F��hZ�����1��7�3�2��C�������
T��_��]���
�8�c�'�0�o�@���P���A�R��U���u�u�u�%�c�����8����U ��h_��F܊� �d�d�
�d�W�W���&ǹ��R
��v'�� ���'�d�
�m�1��B���	���l�N��Uʥ�a��4�0����������@9��P1�Gʢ�0�u�&�9�#�-�(���&����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�b�3��h�O���B�����h=������7�3�0��i�Dց�����9��R�����u�u�u�
��>����0����U��Z��*���
�l�u�=�9�u�����ԓ�V��[�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�c�n�(���H����CU��N������4�0���(����Hǹ��U��_�����h�_�u�u�w�}��������l��@��U¦�9�!�%�'�0�o�C���P���A�R��U���u�u�u�%�c�����8����U ��h_��G���2�c�c�_�w�}�(ہ�����r/��B����
�e�3�
�b�d����D���F�N��A���4�0��
�"�;���&����T9��N�����&�9�!�%�%�:�E��Q���A��N�����u�u�u�u�'�i�$�������Q��R��A��
� �d�f��n�}���Y����`��R
��*���3�'�d�
�f�;�(��O����[�N��U���%�a��4�2��(�������9��E��B��"�0�u�&�;�)�܁�����
U�N��R��u�9�0�_�w�}�W���&ǹ��R
��v'�� ���'�d�
�e�1��B���	��ƹF��hZ�����1��7�3�2��C�������T��N�U���u�u�u�%�c�����8����U ��h_��G���2�c�c�"�2�}��������A��^�]���h�r�r�u�;�8�}���Y���C9��d�����
� �3�'�f��(���H����CU��N������4�0���(����Hǹ��U��\�����h�_�u�u�w�}��������l��@��U¦�9�!�%�
�2��G��I���W����ߊu�u�u�u����������F ��E1�*ߊ�0�
�c�n�w�}����*����W'��U�����a�b�3�
�d�k����D���F�N��A���4�0��
�"�;���&ƹ��T9��N�����&�9�!�%�%�:�E��Q���A��N�����u�u�u�u�'�i�$�������Q��R��A���3�
�f�l�'�f�W���	�ғ�P��S/�����0�
�a�m�1��D���	���l�N��Uʥ�a��4�0����������9��P1�Gʢ�0�u�&�9�#�-�(���&����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�
� �f�n�(��s���C9��d�����
� �3�'�f��G���&����l��S��U���u�u�2�%�1��D߁�Kӑ��]F��R����
�0�
�d�a�m�W���H����_��=N��U���u�
�
�6�;�9�>�������S��h��*��n�u�u�%�c�����8����U ��h_��Dۊ� �d�e�
�d�a�W���Y�����h=������7�3�0��h�N���������YN�����8�d�
�0��l�A��Y���O��[�����u�u�u�
��>����0����U��[��E���
�`�`�%�l�}�WϮ�M����_��~1�����
�`�d�
�"�l�Gց�J���9F�N��U���
�6�9�1��?����&�ӓ�l��hY�U���;�}�0�
�:�l�(���&����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�d�3��k�E���B�����h=������7�3�0��h�F܁�����9��R�����u�u�u�
��>����0����U��[��*���
�e�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���C9��d�����
� �3�'�f��E���&����l��=N��U���
�6�9�1��?����&�ӓ�9��h_�F���u�h�_�u�w�}�W���&����D��F��*���
�%�!�
�2����&����W��h��*���}�|�h�r�p�}����s���F�G1��&���0��
� �1�/�Fځ�O����lQ��d��Uʥ�a��4�0����������^��B1�Fڊ�f�i�u�u�w�}�WϮ�M����_��~1�����
�`�d�
�2��E������R��R	�����
�0�
�8�f�����H�Г�CV��C_��\��r�r�u�9�2�W�W���Y�Ƽ�9��V��4��� �3�'�d��j����O�Փ� ]ǻN��*ފ�6�9�1��5�;����L����U��]�����h�_�u�u�w�}�(ہ�����r/��B����
�c�'�2�`�j� ���Yۇ��A��G�����9�!�%�a�%�:�E��&����Z��G��U��|�0�&�u�w�}�W���	�ғ�P��S/�����0�
�`�d��(�F��&����F�G1��&���0��
� �1�/�Fځ�&����S��G]��H�ߊu�u�u�u�%����I����D��F�����%�l�'�2�e�k�_���D����F��D��U���u�u�%�a��<����&����V��1����f�_�u�u����������F ��E1�*���3�
�c�a�'�}�J�ԜY���F��1������
� �3�%�l�(�������Q��_��]���'�2�%�&�0�.����	�Փ�V��_�����<�d�e�u�w�l�^ϻ�
��ƹF�N��*ފ�6�9�1��5�;����L����U��]����u�u�%�a��<����&����V��1�*���d�`�
�f�k�}�W���Y����lR��T�����7�3�0�
�b�l�(���&����D��F��*���
�%�!�
�2����&����W��h��*���}�|�h�r�p�}����s���F�G1��&���0��
� �1�/�Fځ�I����P��h����u�
�
�6�;�9�>�������S��1��*��m�%�u�h�]�}�W���Y����R��@��U´�
�0�
�%�#���������A��_�*���
�!�}�|�j�z�P������F�N������4�0���(����Hƹ��l��hY�N���u�%�a��6�8�6�������lW��]�� ��c�
�f�i�w�}�W���YӖ��l5��[��<���3�0�
�`�f�����L�ƻ�V�V�����%�!�
�0��0�Fف�����S��G^�����|�h�r�r�w�1��ԜY���F��1������
� �3�%�l�(�������^��UךU���
�
�6�9�3���������lT��Q��C���%�u�h�_�w�}�W���&ǹ��R
��v'�� ���'�d�
�a�%�:�@��������E�����2�&�9�!�'�h����K����C��^�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�b�o�(���H����CU��N������4�0���(����Hƹ��l ��X�*��i�u�u�u�w�}����*����W'��U�����`�d�
�0��h�W����έ�l��h�����0�
�8�d��8�(��O����l��^��H��r�u�9�0�]�}�W���Y����`��R
��*���3�'�d�
�c�;�(��K����9F���*���9�1��7�1�8�(���KŹ��lW��1��U��_�u�u�u�w��(�������l��Q��Dߊ�a�'�2�b�d�*��������T9��D�����!�%�f�'�0�o�Fځ�	ù��N��S��D���0�&�u�u�w�}�WϮ�M����_��~1�����
�`�g�
�"�l�@ց�J���F��1������
� �3�%�l�(�������
U��N�U���u�u�u�%�c�����8����U ��h_��Dފ�0�
�`�u�?�3�_�������C��h��*���d�
�0�
�f�k�������F�_��U���0�_�u�u�w�}�(ہ�����r/��B����
�c�3�
�a�k���Y����lR��T�����7�3�0�
�b�o�(���H����CU�
NךU���u�u�0�
�c�}����Q����V��G��*���
�8�d�
�2��F���	�֓�GW�N��R��u�9�0�_�w�}�W���&ǹ��R
��v'�� ���'�d�
�
�2��@��Y����lR��T�����7�3�0�
�b�o�(���H����CU�
NךU���u�u�
�
�4�1��������A9��h�����b�u�=�;��-����	����l��h��D݊�0�
�d�f�'�m���I���W����ߊu�u�u�u����������F ��E1�*���3�
�b�e�'�f�W���	�ғ�P��S/�����0�
�`�f��(�F��&���FǻN��U���
�
�6�9�3���������l��R	��B���=�;�}�%�%�:��������l��X�����d�`�%�e�>�l�G���Y�����RNךU���u�u�
�
�4�1��������A9��h\�����b�b�%�n�w�}����*����W'��U�����`�f�
� �f�o�(��E��ƹF�N��*ފ�6�9�1��5�;����J����V�� W�����}�%�'�2�'�.��������S��R	��D���%�e�<�d�g�}�W��PӃ��VFǻN��U���
�
�6�9�3���������lU��Q��B���%�n�u�u�'�i�$�������Q��R��@��
� �d�g��n�K���Y���F��hZ�����1��7�3�2��D�������_��_��]���'�2�%�&�0�.����	�ғ�V��\�����<�d�e�u�w�l�^ϻ�
��ƹF�N��*ފ�6�9�1��5�;����L����U�� \����u�u�%�a��<����&����V��1�*���d�f�
�f�k�}�W���Y����lR��T�����7�3�0�
�d�.����N����[�������%�&�2�&�;�)��������W��G����e�u�u�d�~�8����Y���F��hZ�����1��7�3�2��B��&����T��G]�U���%�a��4�2��(�������9��h��D��
�f�i�u�w�}�W���	�ғ�P��S/�����0�
�f�&�%�:�@��������E�����2�&�9�!�'�d����K����C��^�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�b�n�(���H����CU��N������4�0���(����Hƹ��l ��Y�*��i�u�u�u�w�}����*����W'��U�����`�&�'�2�o�h� ���Yۇ��A��G�����9�!�%�m�%�:�E��&����Z��G��U��|�0�&�u�w�}�W�������T��N������4�0���(����Hƹ��l ��Y�*��i�u�u�u�w�}����*����W'��U�����`�&�'�2�o�h� ���Yۇ��A��G�����9�!�%�b�%�:�E��&����Z��G��U��|�0�&�u�w�}�W���	�ғ�P��S/�����0�
�`�f��(�F��&����F�G1��&���0��
� �1�/�Fځ�N����Q��h�I���u�u�u�u�'�i�$�������Q��R��@���'�2�m�`� �8�Wǿ�&����C��P1�����%�c�'�2�e�i�(���&����O�I�\ʰ�&�u�u�u�w�}����*����W'��U�����`�f�
� �f�h�(��s���C9��d�����
� �3�'�f��O���&����l��S��U���u�u�%�a��<����&����V��1�����m�`�"�0�w�<�(���&����T9��[1�����'�2�g�f��-�(���Q���A��N�����u�u�u�u�'�i�$�������Q��R��@��
� �d�c��n�}���Y����`��R
��*���3�'�d�
�n�;�(��N����[�N��U���%�a��4�2��(�������9��E��M���"�0�u�4��8�(�������_9��G_�����g�g�
�%��)�_���D����F��D��U���u�u�%�a��<����&����V��1�*���d�b�
�f�]�}�W���&����V��h�����d�
�
� �f�k�(��E��ƹF�N����� �m�e�%�w�5��������CW��E��G��}�|�h�r�p�}����s���F�G1��&���0��
� �1�/�Fځ�&����R��=N��U���
�6�9�1��?����&�ӓ�9��h_�A���u�h�_�u�w�}�W���&����V��h�����d�
�
�0��m�W����έ�l��h�����0�
�8�d��8�(��L����l��^��H��r�u�9�0�]�}�W���Y����`��R
��*���3�'�d�
�n�;�(��N����9F���*���9�1��7�1�8�(���M¹��lW��1��U��_�u�u�u�w��(�������l��Q��Dߊ�
�0�
�e�w�5����	����l��C	�����8�d�
�0��l�A���I����V�
N��R���9�0�_�u�w�}�W���&����V��h�����d�
�e�3��j�C���B�����h=������7�3�0��h�C���&����l��S��U���u�u�%�a��<����&����V��1�����c�l�"�0�w�.����	�ߓ�V��X�E���u�d�|�0�$�}�W���Y����lR��T�����7�3�0�
�b�n����L�֓� ]ǻN��*ފ�6�9�1��5�;����L�Г�F9�� Z��F��u�u�u�u�w�:����&����CT��_��]���
�8�d�
�2��F��I���W����ߊu�u�u�u����������F ��E1�*ߊ�0�
�b�n�w�}����*����W'��U�����`�b�3�
�b�l����D���F�N��A���4�0��
�"�;���&ƹ��T9��N�����&�9�!�%�d�/���H����[�I�����u�u�u�u�w�-�C�������z9��Q��*���c�3�
�`�c�-�L���YӖ��l5��[��<���3�0�
�`�o�;�(��A����[�N��U���%�a��4�2��(�������9��E��C���"�0�u�&�;�)��������P��G��U��|�0�&�u�w�}�W���	�ғ�P��S/�����0�
�`�b�1��B���	��ƓF�C��*݊�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(߁�	����l��D�����2�
�'�6�m�-����
ۖ��l$��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b��e�4��1�^������F�N��U���%�b��e�6���������Z�G1��7���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*ڊ�;�&�2�4�$�:�W�������K��N������e�<�
�>���������PF��G�����%�b��e�w��(���&����F�� 1��E���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��9��h��\���=�;�_�u�w�}�W���Y����q9��^ �����h�%�b��g�W�W���Y�Ʃ�@�N��U���u�u�%�b��m���������h,��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����l��A�����<�u�&�<�9�-����
���9F���*���e�4�
�9��3��������]9��X��U���6�&�}�
���G���&������h,��E���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lQ��h_�����9�|�u�=�9�W�W���Y���F�� 1��Dڊ�%�#�1�<��4�W��	�ѓ�lW��V����u�u�u�u�2�.�W���Y���F���*���e�4�
�9��3����E�Ƽ�9��^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l$��1��*���u�&�<�;�'�2����Y��ƹF��hY��*���<�
�<�
�$�4��������C��R������d�y�%�`��F߁����C9��u1�*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�N����9��h��\���=�;�_�u�w�}�W���Y����q9��h�����i�u�
�
��m�}���Y���V
��d��U���u�u�u�%�`��F߁�����Z�G1��7��
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����q9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�d�4��1�(���
����@��Y1�����u�'�6�&���(���H����E
����*���d�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*���4�
�9�|�w�5��ԜY���F�N��B���d�
�%�#�3�4�(���Y����lQ��h_�����9�n�u�u�w�}����Y���F�N��U���
�
�d�4��1�(���
���F�� 1��Dۊ�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h,��D���
�<�u�&�>�3�������KǻN��*݊�
�d�<�
�>���������PF��G�����%�b��d�{�-�@���H¹��V�G1��7��
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l$��1��*���|�u�=�;�]�}�W���Y���C9��u1�*���&�2�i�u���(��s���F�R��U���u�u�u�u�w�-�@���H¹��l��R������d�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��u1�*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
�e�<�(���&����Z��D�����:�u�u�'�4�.�_���&����l��A��U���
�
�g�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�
�g�4�
�;�t�W������F�N��Uʥ�b��d�
�'�+����&����[��hY��*���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
�e�<�(���&����Z�
N��B���d�
�%�#�3�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���g�<�
�<�w�.����	����@�CךU���
�
�
�g�>�����
����l��TN����0�&�%�b��l�[Ϯ�N����9��R	�����d�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h,��G���
�9�|�u�?�3�}���Y���F�G1��7��
�;�&�2�k�}�(؁�&����F�N�����u�u�u�u�w�}�WϮ�N����9��h��U��%�b��d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��7��
�%�#�1�>�����
������T��[���_�u�u�
���D���&����Z��^	�����;�%�:�u�w�/����Q����q9��h�����u�
�
�
�d�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�f�6�����Y����l�N��U���u�%�b��f���������@��S��*݊�
�f�4�
�;�f�W���Y����_��=N��U���u�u�u�
���D���&����Z��^	��Hʥ�b��d�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�f�<��4�W�������A	��D�X�ߊu�u�
�
��n��������@��h����%�:�0�&�'�j�5��UӖ��l$��1�����%�b��d��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���f�4�
�9�~�}����s���F�N������d�
�;�$�:�K���&Ĺ��U��N��U���0�&�u�u�w�}�W���YӖ��l$��1��*���u�h�%�b��l�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����d�
�%�!�9�����ƭ�@�������{�x�_�u�w��(���M����E
��^ �����&�<�;�%�8�}�W�������C9��u1�*���#�1�u�
���C���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��i�������G��d��U���u�u�u�%�`��Fہ�	����l��D��I���
�
�
�a�6����Y���F��[�����u�u�u�u�w��(���M����E
��^ �����h�%�b��f���������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
�c�4�(���Y����T��E�����x�_�u�u���(�������T9��D��*���6�o�%�:�2�.����;������h,��A���0�y�%�b��l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�a�4��1�^������F�N��U���%�b��d��3����E�Ƽ�9��Z�U���u�u�0�&�w�}�W���Y�����h,��A���
�<�u�h�'�j�5��&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b��d��-��������TF��D��U���6�&�{�x�]�}�W���&����l��A�����<�
�&�<�9�-����Y����V��G1��7��
�%�#�1�w��(���L����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(�������WO�C��U���u�u�u�u�w�-�@���Hƹ��l��h�����i�u�
�
��h������ƹF�N�����_�u�u�u�w�}�W���&����l��A�����<�u�h�%�`��Fځ�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
���B���&����R��P �����&�{�x�_�w�}�(؁�&�ӓ�]9��P1�����
�'�6�o�'�2����	�ѓ�lW����*���`�%�0�y�'�j�5��&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�b�<�(���P�Ƹ�V�N��U���u�u�%�b��l�(���
���F�� 1��D��u�u�u�u�2�.�W���Y���F���*���`�<�
�<�w�`����;����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b��l��������l�������%�:�0�&�w�p�W���	�ѓ�lW��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��B���d�4�
�9�{�-�@���H����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(ށ�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�@���H����E
��^ �����h�%�b��f�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b��d�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l$��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��*ۊ�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(؁�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�b��d�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h,��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.����;�ԓ�C9��SB��*݊�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��7���4�
�9�|�w�5��ԜY���F�N��B���g�4�
�9��3����E�Ƽ�9��1��*���n�u�u�u�w�8����Y���F�N��*݊�
�
�%�#�3�4�(���Y����lQ��h\�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l$��h�����4�&�2�u�%�>���T���F�� 1��G���
�<�
�&�>�3����Y�Ƽ�\��DF��B���g�u�
�
������Y����q9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(؁�&����l��R������g�_�u�w�}�W������F�N��Uʥ�b��g�<��4�W��	�ѓ�lT��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(܁�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��1��*���
�;�&�2�6�.���������T��]���
�
�
�%�!�9�W���&����R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@���J����E
��N�����u�u�u�u�w�}����;�Փ�C9��S1��*���u�h�%�b��n������ƹF�N�����_�u�u�u�w�}�W���&����R��[
�����2�i�u�
���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
������Ӈ��Z��G�����u�x�u�u�'�j�5�������T9��D��*���6�o�%�:�2�.����;���C9��u1�����y�%�b��d�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��B���f�4�
�9�~�}����s���F�N������f�<�
�>�}�JϮ�N����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lU��Y1����u�
�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��7���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�b��i��������l��h�����%�:�u�u�%�>����&Ĺ��9��h��Yʥ�b��a�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�
�
�%�#�3�t����Y���F�N��U���
�
�
�%�!�9���������h,��*���#�1�_�u�w�}�W������F�N��Uʥ�b��a�4��1�(���
���F�� 1��A���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��u1�����<�u�&�<�9�-����
���9F���*���
�;�&�2�6�.���������T��]���
�
�y�%�`��C�������lQ��hZ�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����;�ғ�C9��SG�����u�u�u�u�w�}�WϮ�N����l��D��I���
�
�
�n�w�}�W�������9F�N��U���u�
�
�
��3����E�Ƽ�9��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@���L����E
��^ �����&�<�;�%�8�8����T�����h,��*���#�1�<�
�>���������PF��G�����%�b��`�6����	�ѓ�lS��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&Ĺ��9��h��*���&�2�i�u���(ځ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�lS��G1�����
�<�u�h�'�j�5�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`��B���&����R��P �����&�{�x�_�w�}�(؁�&ƹ��l��h�����%�:�u�u�%�>����&Ĺ��J��hY��*ߊ�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����q9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��1��*���u�h�%�b��h����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(ف�	����l��D�����2�
�'�6�m�-����
ۖ��l$��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b��c�4��1�^������F�N��U���%�b��c�6���������Z�G1��7���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*܊�;�&�2�4�$�:�W�������K��N������c�<�
�>���������PF��G�����%�b��c�w��(���&����F�� 1��C���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��9��h��\���=�;�_�u�w�}�W���Y����q9��^ �����h�%�b��a�W�W���Y�Ʃ�@�N��U���u�u�%�b��k���������h,��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1��7���4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�9�� 1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ѓ�lQ��G1�����!�0�u�u�w�}�W���YӖ��l$��h�����<�
�<�u�j�-�@���N����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9�� 1��*���
�;�&�2�k�}�(؁�&Ĺ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�N����l��D�����2�
�'�6�m�-����
ۖ��l$��N��B���b�%�0�y�'�j�5�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b��b�6�����Y����l�N��U���u�%�b��`�4�(���Y����lQ��hY�U���u�u�0�&�w�}�W���Y�����h,��*���&�2�i�u���(؁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b��m�4��1�(���
����@��YN�����&�u�x�u�w�-�@���A����E
��^ �����&�<�;�%�8�}�W�������C9��u1�����9�y�%�b��e��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*݊�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�b��e��������l��R������m�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���m�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q����;�ޓ�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l$��h�����|�!�0�u�w�}�W���Y����lQ��hV�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ׁ�����Z�G1��7���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�l_��G1�����
�<�u�&�>�3�������KǻN��*݊�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�`��N���&������h,��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��1��*���|�u�=�;�]�}�W���Y���C9��u1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h,��*���#�1�<�
�>�}�JϮ�N����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����;�ߓ�]9��PN�����u�'�6�&�y�p�}���Y����q9��^ �����&�<�;�%�8�}�W�������C9��u1�U���
�
�
�'�0�}�(؁�&ʹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F�� 1��L�ߊu�u�u�u�;�8�}���Y���F�G1��7���<�
�<�u�j�-�@���@����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hW��*ڊ�%�#�1�u���(߁�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l��m�������G��d��U���u�u�u�%�n��G���&����Z��^	��Hʥ�l��e�4��1�L���Y�����RNךU���u�u�u�u���(߁�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�l��g�4�(���&����T��E��Oʥ�:�0�&�%�n��G���&ʹ��9��R	�����e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��z1�����9�|�u�=�9�W�W���Y���F��1��E���
�<�u�h�'�d�:��s���F�R��U���u�u�u�u�w�-�N���I����@��S��*ӊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��^�����1�<�
�<�w�.����	����@�CךU���
�
�
�e�6���������l��^	�����u�u�'�6�$�u�(ց�&�֓�C9��SB��*ӊ�
�e�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���e�4�
�9�~�}����s���F�N������d�
�%�!�9���������h#��E���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�e�6���������Z�G1��8��
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hW��*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�e�<��4�(�������A	��N�����&�%�l��f�q����4����C��N��L���d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����l_��h_�����9�|�u�=�9�W�W���Y���F��1��Dڊ�;�&�2�i�w��(���I���F�N�����u�u�u�u�w�}����4����Z��^	��Hʥ�l��d�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1��Dۊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��l��������l��h�����%�:�u�u�%�>����&ʹ��W��G1�����
�
�
�d�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�d�4��1�^������F�N��U���%�l��d��-��������TF���*���d�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
��l��������l��R������d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ӊ�
�d�<�
�>�}����Ӗ��P��N����u�
�
�
�f�4�(���&����T��E��Oʥ�:�0�&�%�n��F��	�ߓ�lW��G��Yʥ�l��d�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hW��*���4�
�9�|�w�5��ԜY���F�N��L���d�
�;�&�0�a�W���&����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�lW��^ �����h�%�l��f�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��L���d�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(�������W9��h��*���<�;�%�:�w�}����
�μ�
9��\�����1�u�
�
��o��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�e�<�(���P�Ƹ�V�N��U���u�u�%�l��l�(�������]9��PN�U���
�
�g�4��1�L���Y�����RNךU���u�u�u�u���(�������W9��h��U��%�l��d��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�
�g�>�����
������T��[���_�u�u�
���E���&����R��P �����o�%�:�0�$�-�N���H����l_��h_�����y�%�l��f��������F��P��U���u�u�<�u��-��������Z��S��*ӊ�
�g�4�
�;�t�W������F�N��Uʥ�l��d�
�9�.���Y����~9��d��U���u�0�&�u�w�}�W���Y����l_��h_�����<�u�h�%�n��F݁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�l��d�
�'�+����&����R��P �����&�{�x�_�w�}�(ց�&�Փ�C9��S1��*���
�&�<�;�'�2�W�������@N��1��Dي�%�#�1�u���(�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
���D���&����F��R ��U���u�u�u�u�'�d�:��&����_��Y1����u�
�
�
�d�<�(���B���F����ߊu�u�u�u�w�}�(ց�&�Փ�C9��S1��*���u�h�%�l��l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
��n�����ƭ�@�������{�x�_�u�w��(���J����@��V�����'�6�o�%�8�8�Ǯ�@���� J��hW��*���%�0�y�%�n��F܁�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�f�6�����Y����l�N��U���u�%�l��f��������C9��z1�N���u�u�u�0�$�}�W���Y���F��hW��*���<�
�<�u�j�-�N���H����V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�l��f���������@��V�����'�6�&�{�z�W�W���&ʹ��R��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��L���d�
�%�#�3�}�(ց�&�ғ�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���M����E
��N�����u�u�u�u�w�}����4����R��[
�����2�i�u�
���C���&����9F�N��U���0�_�u�u�w�}�W���&ʹ��R��G1�����
�<�u�h�'�d�:��&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(�������TF��D��U���6�&�{�x�]�}�W���&����l��D�����2�
�'�6�m�-����
ۖ��l+��B��*ӊ�
�a�%�0�{�-�N���Hǹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
��i�������G��d��U���u�u�u�%�n��Fہ�����Z�G1��8��n�u�u�u�w�8����Y���F�N��*ӊ�
�a�<�
�>�}�JϮ�@����9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n��Fځ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��[�����1�<�
�<��.����	����	F��X��¥�l��d�
�'�+����&ʹ��S��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����l��A��\ʡ�0�u�u�u�w�}�W���	�ߓ�lW��V�����;�&�2�i�w��(���L����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�
9��[�����1�<�
�<�w�`����4����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ց�&�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����~9��h�����4�&�2�
�%�>�MϮ�������h#��@���
�
�
�`�'�8�[Ϯ�@����9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(�������WO�C��U���u�u�u�u�w�-�N���Hƹ��l��R������d�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�`�>�����DӖ��l+��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�N���H����E
��^ �����&�<�;�%�8�8����T�����h#��*���#�1�<�
�>���������PF��G�����%�l��d�6����	�ߓ�lW��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&ʹ��9��h��*���&�2�i�u���(ށ�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�lW��G1�����
�<�u�h�'�d�:�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n��F���&����R��P �����&�{�x�_�w�}�(ց�&¹��l��h�����%�:�u�u�%�>����&ʹ��J��hW��*ۊ�'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����~9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�
9��1��*���u�h�%�l��l����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ӊ�
�
�%�#�3�4�(���Y����T��E�����x�_�u�u���(݁�	����l��D�����2�
�'�6�m�-����
ۖ��l+��h�����u�
�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�l��g�4��1�^������F�N��U���%�l��g�6���������Z�G1��8���4�
�9�n�w�}�W�������9F�N��U���u�
�
�
��-��������TF���*���
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hW��*؊�;�&�2�4�$�:�W�������K��N������g�<�
�>���������PF��G�����%�l��g�w��(���&����F��1��G���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ʹ��9��h��\���=�;�_�u�w�}�W���Y����~9��^ �����h�%�l��e�W�W���Y�Ʃ�@�N��U���u�u�%�l��o���������h#��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R��[
�����2�4�&�2�w�/����W���F�G1��8���4�
�9�
�9�.����
����C��T�����&�}�
�
�������Ƽ�
9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ߓ�lU��G1�����!�0�u�u�w�}�W���YӖ��l+��h�����<�
�<�u�j�-�N���J����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�
9��1��*���
�;�&�2�k�}�(ց�&����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�@����l��D�����2�
�'�6�m�-����
ۖ��l+��N��L���f�%�0�y�'�d�:�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�l��f�6�����Y����l�N��U���u�%�l��d�4�(���Y����l_��h]�U���u�u�0�&�w�}�W���Y�����h#��*���&�2�i�u���(܁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�l��a�4��1�(���
����@��YN�����&�u�x�u�w�-�N���M����E
��^ �����&�<�;�%�8�}�W�������C9��z1�����9�y�%�l��i��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
��-����PӒ��]FǻN��U���u�u�
�
����������@��S��*ӊ�
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�l��i��������l��R������a�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��L���a�<�
�<�w�.����	����@�CךU���
�
�
�
�9�.����
����C��T�����&�}�
�
��q����4�ғ�A����*���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l+��h�����|�!�0�u�w�}�W���Y����l_��hZ�����2�i�u�
���L���Y�����RNךU���u�u�u�u���(ہ�����Z�G1��8���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�lS��G1�����
�<�u�&�>�3�������KǻN��*ӊ�
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�n��B���&������h#��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�
9��1��*���|�u�=�;�]�}�W���Y���C9��z1�����9�
�;�&�0�a�W���&����R��[
�U���u�u�0�&�w�}�W���Y�����h#��*���#�1�<�
�>�}�JϮ�@����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����4�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����~9��^ �����&�<�;�%�8�}�W�������C9��z1�U���
�
�
�'�0�}�(ց�&ƹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
����������[��=N��U���u�u�u�
���(���
���F��1��@�ߊu�u�u�u�;�8�}���Y���F�G1��8���<�
�<�u�j�-�N���L����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����R��[
�����2�4�&�2��/���	����@��hW��*܊�%�#�1�u���(ف�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l��k�������G��d��U���u�u�u�%�n��A���&����Z��^	��Hʥ�l��c�4��1�L���Y�����RNךU���u�u�u�u���(ف�	����l��D��I���
�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�l��a�4�(���&����T��E��Oʥ�:�0�&�%�n��A���&ʹ��9��R	�����c�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��z1�����9�|�u�=�9�W�W���Y���F��1��C���
�<�u�h�'�d�:��s���F�R��U���u�u�u�u�w�-�N���O����@��S��*ӊ�
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9�� 1��*���
�;�&�2�6�.��������@H�d��Uʥ�l��b�4��1�(���
����@��Y1�����u�'�6�&���(���&����_�G1��8���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h#��*���#�1�|�!�2�}�W���Y���F��hW��*݊�%�#�1�<��4�W��	�ߓ�lQ��G1���ߊu�u�u�u�;�8�}���Y���F�G1��8���4�
�9�
�9�.���Y����~9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ʹ��9��h��U���<�;�%�:�2�.�W��Y����l_��hY�����2�4�&�2��/���	����@��hW��*���%�l��b�'�8�[Ϯ�@����l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�n��@���&����F��R ��U���u�u�u�u�'�d�:�������TF���*���n�u�u�u�w�8����Y���F�N��*ӊ�
�
�;�&�0�a�W���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�l��e��������l�������%�:�0�&�w�p�W���	�ߓ�l^��G1�����
�<�
�&�>�3����Y�Ƽ�\��DF��L���m�4�
�9�{�-�N���A����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(ׁ�	����O��_�����u�u�u�u�w��(���&����_��Y1����u�
�
�
��-����s���F�R��U���u�u�u�u�w�-�N���A����E
��^ �����h�%�l��o�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�l��m�>�����
������T��[���_�u�u�
���(���
����@��Y1�����u�'�6�&���(���UӖ��l+��h�����
�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hW��*Ҋ�%�#�1�|�#�8�W���Y���F���*���
�;�&�2�k�}�(ց�&��ƹF�N�����_�u�u�u�w�}�W���&����Z��^	��Hʥ�l��m�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h#��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�
��-��������T9��D��*���6�o�%�:�2�.����4�ߓ�C9��SB��*ӊ�
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��8���4�
�9�|�w�5��ԜY���F�N��L���l�4�
�9��3����E�Ƽ�
9��1��*���n�u�u�u�w�8����Y���F�N��*ӊ�
�
�%�#�3�4�(���Y����l_��hW�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l+��h�����4�&�2�u�%�>���T���F��1��L���
�<�
�&�>�3����Y�Ƽ�\��DF��L���l�u�
�
������Y����~9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(ց�&ʹ��l��R������l�_�u�w�}�W������F�N��Uʥ�l��l�<��4�W��	�ߓ�l_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�0�
�:�l�(���H����CU�
NךU���u�u�
�
������ӑ��]F��R�����3�
�b�
�e�m�W���H����_��=N��U���u�0�
�8�n�;�(��H����9F���*���d�
� �d�c��D��Y���F���*���e�<�
�<�w�5��������C^��B1�E���}�|�h�r�p�}����s���F�D�����e�3�
�e�o�-�L���Yӕ��l��\�� ��`�
�f�i�w�}�W���YӖ��l+��1��*���u�=�;�}�2���������9��^��H��r�u�9�0�]�}�W���Y����G��1��*��`�%�n�u�w�.����	�Փ�F9�� V��G��u�d�u�=�9�u�;���&����	��h[��*��
�
� �d�`��E������]��[��F���9�0�w�w�]�}�W���&����9��h_�A���u�h�w�w� �8�WǷ�&����\��X��@���e�e�!�3��m�E���Y�ƭ�l��D��ފ�|�0�&�u�g�f�W���
����^��h��D��
�g�i�u�f�}����Q����Z9��E1�����
�
�g�
��(�F��&�����T�����a�b�u�9�2��U�ԜY�ƿ�_9��G_�����e�c�%�u�j��Uϩ�����9��h(��*���%�`�d�e�g�)����I�ԓ�F�V�����
�#�
�|�2�.�W��B�����h��D݊� �d�e�
�e�a�W��Y����N��h��3����:�
�
��o�(�������9��S�����;�!�9�a��}����[����F�D�����m�3�
�d�o�-�W��[����[�������:�
�:�%�b�l�G�������V��h�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����8�d�
� �f�l�(��E���F��R �����<��'��8��(ށ�Kù��U��Y�����u�%�6�;�#�1�C��Y����D��d��Uʦ�9�!�%�
�"�e�A���Y���D��_��]���
� �m�g�'�}�W�������l
��h-�����u�e�n�u�w�.����	�֓�F9��^��F��u�u�u�u�w�-�N���J����@��@��U¦�9�!�%�f�1��G���	����[�I�����u�u�u�u�w�-�N���Hƹ��l��d��Uʦ�9�!�%�d�1��E���	���l�N��Uʥ�l��`�<��4�W����ο�_9��G_�����e�a�%�}�~�`�P���Y����l�N��Uʦ�9�!�%�e�1��E���	��ƹF��R����
� �d�`��n�K���Y���F��hW��*݊�;�&�2�"�2�}��������l ��^�*��e�u�u�d�~�8����Y���F��R����
� �d�a��n�}���Y����G��1��*��e�%�u�h�]�}�W���Y����~9��^ �����=�;�}�0��0�Fف�����9��^��H��r�u�9�0�]�}�W���Y����G��1��*��f�%�n�u�w�.����	�ғ�F9��Y��F��u�u�u�u�w�-�N���H¹��l�������0�
�8�d��(�F��&���F�_��U���0�_�u�u�w�}��������U��X����u�u�&�9�#�-�B���&����l��S��U���u�u�%�l��l�(���
����[����*���d�
� �d�g��E��Y���O��[�����u�u�u�0��0�Eہ�����9��d��Uʦ�9�!�%�
�"�e�E���Y���D��_��]���
� �m�g�'�}�W�������l
��hZ�����u�e�n�u�w�.����	����l^��h�I���d�u�=�;��0�(���A�ԓ�F�V�����
�#�
�|�2�.�W��B�����h��A���
�c�
�g�k�}�F������G��Q��@؊�d�h�4�
�8�.�(���&����_��^�����u�0�
�8�b�;�(��A����[�N��U���%�l��g�>��������@��C�����`�
�g�e�w�}�F�������9F�N��U���
�
�a�<��4�L���Yӕ��l��1��*��
�g�i�u�f�}����Q����U��\��D��4�
�:�&��+�(�������V�=N��U���
�8�b�3��m�C���Y���F�N������a�<�
�>�}����Q����G��h��M���%�}�|�h�p�z�W������F�N�����%�
� �d�f��D�ԜY�ƿ�_9��GV�� ��e�%�u�h�u�� ���Yے��l ��[�����u�%�6�;�#�1�C���Y����D��d��Uʦ�9�!�%�
�"�l�Dށ�J���9F�N��U���
�
�
�;�$�:� ���Yە��l��1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�b�3�
�g�i���Y����V
��Z�� ��c�%�u�h�u�� ���Yے��l ��[�����u�%�6�;�#�1�C��Y����D��d��Uʡ�%�3�
�`��l�K���5����u	��{��*ߊ�=�
� �m�e�-�_���Y�ƨ�D��^����u�0�4�n�