-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�m�l��m��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e� �&�4�2��(���Y����g"��x)��*�����}�`�3�*����P���F��h��Oʜ�u��
���f�W���	�֓�]��[��<���4�
�9�u�w��$���5����l�N��E���&�4�0���}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��D�����
�
�%�#�3�g�>���-����t/��=N��U���
�;�6�9�3��E��0�Ɵ�w9��p'��#����u�d�u�8�3���B�����h;�����1��g�4��1�W���7ӵ��l*��~-�U���%�e� �&�6�8�6���Y�ƅ�5��h"��<������}�b�9� ���Y����F�G1�� ���4�0��
��-����Cӯ��`2��{!��6�ߊu�u�
�
�9�>����0���/��d:��9�������w�l�W������]ǻN��*ڊ�;�6�9�1��i��������z(��c*��:���n�u�u�%�g���������F��~ ��!�����
����_������\F��d��Uʥ�e� �&�4�2��(ځ�	����\��yN��1�����_�u�w��(�������r/��T��;ʆ�������8���H�ƨ�D��^����u�
�
�;�4�1����O����E
��N��U���
���n�w�}����,����_��~1�Oʜ�u��
����2���+������Y��E��u�u�%�e��.����8����R��[
��U��������W�W���&ù��@��R
��*���u������4���:����W��S�����|�_�u�u����������l^��G1�����u��
���L���YӖ��l3��T�����l�o��u���8���&����|4�[�����:�e�n�u�w�-�G���
����W'��1��*���u�u�����0���s���C9��b ������
�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I����P��S/��Dڊ�%�#�1�o��}�#���6����9F���*���6�9�1��f�}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��D�����
�d�4�
�;�}�W���*����|!��d��Uʥ�e� �&�4�2��(��Cӯ��`2��{!��6�����u�d�w�2����I��ƹF��h^�����9�1��d��-����Cӯ��`2��{!��6�ߊu�u�
�
�9�>����0����	F��=��*����
����u�BϺ�����O��N����� �&�4�0���D���&����	F��=��*����n�u�u�'�m�"�������z9��T��;ʆ�������8���H�ƨ�D��^����u�
�
�;�4�1����Hǹ��l��T��;ʆ�����]�}�W���&����R
��v'��@���u��
���(���-���S��X����n�u�u�%�g���������S��G1�����u��
���L���YӖ��l*��^�����0�u�u����;���:����g)��_����!�u�|�_�w�}�(ށ�����v��[�����9�u�u����;���:���F��1�����8�!�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�L����[*��^��*���#�1�o��w�	�(���0��ƹF��h[�����<�<�
�u�w��$���5����l0��c!��]���1�"�!�u�~�W�W���&ƹ��T��Z��D���
�9�u�u���3���>����F�G1��=����8�!�g�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ӓ�Z��^��*؊�%�#�1�o��}�#���6����9F���*���=�<�<�
�w�}�9ύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����{��{�����4�
�9�u�w��$���5����l�N��@���2��8�!�c�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӖ��l.��_"�����
�%�#�1�m��W���&����p]ǻN��*ߊ�<�=�<�<��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��P�����`�4�
�9�w�}�9ύ�=����z%��N������2��8�#�k�Mϗ�Y����)��t1��6���u�d�u�:�9�2�G��Y����lS��^	�����
�
�%�#�3�g�>���-����t/��=N��U���
�<�=�<�>��W���7ӵ��l*��~-��0����}�`�1� �)�W���s���C9����9���!�b�4�
�;�}�W���*����|!��d��Uʥ�`��2��:�)�O��0�Ɵ�w9��p'��#����u�d�u�8�3���B�����h&�����<�
�
�%�!�9�Mϗ�Y����)��tUךU���
�
�<�=�>�4�(���Y����g"��x)��*�����}�`�3�*����P���F��1�����8�!�l�4��1�W���7ӵ��l*��~-�U���%�`��2��0���Y�ƅ�5��h"��<������}�b�9� ���Y����F�G1��=����8�!�d��-����Cӯ��`2��{!��6�ߊu�u�
�
�>�5����&���/��d:��9�������w�l�W������]ǻN��*ߊ�<�=�<�<��l��������z(��c*��:���n�u�u�%�b���������F��~ ��!�����
����_������\F��d��Uʥ�`��2��:�)�F݁�	����\��yN��1�����_�u�w��(�������G9��T��;ʆ�������8���H�ƨ�D��^����u�
�
�<�?�4����J����E
��N��U���
���n�w�}����1����Z��h_�Oʜ�u��
����2���+������Y��E��u�u�%�`��:�;�������R��[
��U��������W�W���&ƹ��T��Z��D���u������4���:����W��S�����|�_�u�u����������S��G1�����u��
���L���YӖ��l*��{����o��u����>���<����N��
�����e�n�u�u�'�j�;�������9��h��U���������}���Y����	��^��*���u������4���:����W��S�����|�_�u�u����������l��A��Oʜ�u��
���f�W���	�ѓ�\��Z��G���u��
���(���-���S��X����n�u�u�%�`�� �������R��[
��U��������W�W���&Ĺ��D*��^��U���������!���6���F��@ ��U���_�u�u�
��2�;����Փ�C9��SN�<����
���l�}�WϮ�N������C1�Oʜ�u��
����2���+������Y��E��u�u�%�b��*����&ǹ��l��T��;ʆ�����]�}�W���&����Z��h[��U���������4���Y����W	��C��\�ߊu�u�
�
�8�����L����E
��N��U���
���n�w�}����5����^��N�<����
�����#���Q����\��XN�N���u�%�b�� �4����&����_�'��&������_�w�}�(؁�����Z��T��;ʆ�������8���H�ƨ�D��^����u�
�
�:��0��������WF��~ ��!�����n�u�w�-�@�������G9��N��U���
���
��	�%���Lӂ��]��G�U���%�b��"�>�4�(ׁ�	����\��yN��1�����_�u�w��(���5����l_�'��&���������W��Y����G	�UךU���
�
�:��:�)�N���&����	F��=��*����n�u�u�'�j�;�������V�'��&���������W��Y����G	�UךU���
�
�:��:�)�F߁�	����\��yN��1�����_�u�w��(���5����lW��N��U���
���
��	�%���Lӂ��]��G�U���%�b��"�>�4�(�������WF��~ ��!�����n�u�w�-�@�������G9��T��;ʆ�������8���H�ƨ�D��^����u�
�
�:��0���&����_�'��&������_�w�}�(؁�����Z��N�<����
�����#���Q����\��XN�N���u�%�b�� �4����J����E
��N��U���
���n�w�}����5����^��Z��U���������4���Y����W	��C��\�ߊu�u�
�
�8�����Hǹ��l��T��;ʆ�����]�}�W���&����Z��h_�Oʜ�u��
����2���+������Y��E��u�u�%�b��*����&�ӓ�C9��SN�<����
���l�}�WϮ�A����Z��V����������4�ԜY�Ƽ�9��Z�����0�
�%�#�3�g�8���*����|!��d��Uʥ�l� �&�4�2���������\��yN��1��������}�F�������V�=N��U���
�;�6�9�3�4��������R��[
��U��������W�W���&�֓�]��[������2��!�m��#ύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����l3��T�����<��2��#�<�(���Y�ƃ�gF��s1��2���_�u�u�
�f���������Z��@'��Oʜ�u��
����2���+������Y��E��u�u�%�d��3��������G*��~ �����1�o��u���8���B�����1�����<�<�u�u���3���>����F�G1�*���4��8�!�6�����Y����g"��x)��N���u�%�d�
�9�>��������\��CN�:���������4���Y����W	��C��\�ߊu�u�
�`��.����5����	��B�����1�o�����;���:����V��=d�����!�6� �0�5�5�ϱ�Y����
P����U���_�u�u�!�%�?����6����v(��v:��;����u�u����}���Y����Z��RN��'���������1���ӄ��R������6� �0�<�]�}�Wͳ�A����^��B�����
�e�a�a�,��(���,����c#��O��9���� �
���`�[���&����g9��o+��EƝ�������J�������_��C�=���������E���I����.��h'�� �����:�=�%�q�;��� ����|%�� @�L��y��
����J��1����j(��g:�����������GÖ�*����l"��
^��9����
��l�`��$���7����W�������u�:�&�4�#�<�(���
����T��N�&������o�w�l�L���YӅ��@��CN��*���&�
�:�<��}�W���&����pF��I�N���u�6�;�!�9�}����&����U��N�&���������W������\F��T��W��n�u�u�6�9�)����	����@��Q��D��������4���Y����\��XN�U��w�e�n�u�w�>�����ƭ�l��D�����e�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�d�l�}�WϽ�����GF��h�����#�c�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���6�;�!�;�w�-��������lV�=��*����
����u�W������F��L�N���u�6�;�!�9�}��������EU��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�D��u�u�6�;�#�3�W�������l
��h^��U���
���
��	�%���Y����G	�N�U��e�e�n�u�w�>�����ƭ�l��D��ފ�u�u��
���(���-��� F��@ ��U���o�u�e�e�u�W�W�������]��G1�����9�a�g�o���;���:����g)��]�����:�e�u�h�u�m�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��H����F�T�����u�%�6�;�#�1�C��Cӵ��l*��~-��0����}�u�:�9�2�G���D����V�=N��U���&�4�!�4��2����ǹ��	F��s1��2������u�d�9� ���Y���F�^�N���u�6�;�!�9�}��������ER��T��!�����
����_�������V�S��E��w�_�u�u�8�.��������]��[��B��������4���Y����\��XN�U��w�d�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�d�g��}���Y����G�������!�9�a�l�m��3���>����v%��eN��U���;�:�e�u�j��G��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���f�1�"�!�w�t�M���H����l�N�����;�u�%�6�9�)����;����g"��x)��*�����}�u�8�3���Y���V��UךU���:�&�4�!�6�����&����pF��d:��9�������w�n��������\�_�E��u�u�6�;�#�3�W�������l
��h*��U���
���
��	�%���Y����G	�N�U��e�w�_�u�w�2����Ӈ��P	��C1��A���o������!���6�����Y��E���h�w�d�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��vN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��_�E��u�u�6�;�#�3�W�������l
��1��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��6��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�4�3����Y����\��h��G���o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�d�n�u�w�>�����ƭ�l��D������o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�d�e�n�w�}��������R��X ��*���g��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�d�d�l�}�WϽ�����GF��h�����#�
�e�o���;���:����g)��Z�����:�e�u�h�u�m�G���s���P	��C��U���6�;�!�9�b�l�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����lǻN�����9�4�
��1�0�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���H��ƹF��C�����u�&�
�;�8�4���
����T]ǻN�����7�!�u�&��3����Ӊ��R��d1����&�2�4�u�$�����B�����Y�����<�
�&�$���ށ�
����	F��s1��2���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:����&ù��@��R
��*ڊ�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��l3��T�����e�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�m�"�������z9��V�����;�&�2�o���;���:���F��P ��U���
�;�6�9�3��G���&����C��T��!�����u�h�p�z�}���Y����R
��h^�����9�1��d�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��E���&�4�0�������Cӵ��l*��~-��0����}�`�1� �)�W���C���V��^�E��e�e�n�u�w�.����Y����f��V��4���
�%�#�1�>�����Y����)��tUךU���<�;�9�%�g���������9��h��*���2�o�����4��Y���9F������%�e� �&�6�8�6���&����Z�=��*����
����u�BϺ�����O��N�����4�u�
�
�9�>����0�ԓ�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*���6�9�1��e�<�(���&����Z�=��*����n�u�u�$�:����&ù��@��R
��*؊�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������r/��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����,����_��~1�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�e� �$�<����&����l��h�����o������}���Y����R
��h^�����9�1��f�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l3��T�����a�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��b ������
�
�'�0�g�$���5����l0��c!��]���1�"�!�u�~�g�W��I����V��^�E��u�u�&�2�6�}�(߁�����V��hZ�����1�<�
�<�w�}�#���6����9F������%�e� �&�6�8�6���&����_��E��Oʆ�����m�}�G��Y����Z��[N��E���&�4�0�����������g"��x)��*�����}�`�3�*����P���F��P ��U���
�;�6�9�3��B�������`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�w�]�}�W�������lV��Y������`�4�
�;���������g"��x)��N���u�&�2�4�w��(�������r/��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�9�>����0�Г�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�g���������9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y����� �&�4�0���(�������]9��PN�&������_�w�}����Ӗ��l3��T�����c�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����,����_��~1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ù��@��R
��*݊�'�2�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��d��Uʦ�2�4�u�
��3��������l��A�����<�u�u����>��Y����Z��[N��E���&�4�0�����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��b ������
�
�;�$�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��h^�����9�1��m�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�I����P��S/��M���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�9�>����0�ޓ�C9��S1�����u��
���}�J���^���F��P ��U���
�;�6�9�3��N���&����	F��s1��2������u�f�}�������9F������%�e� �&�6�8�6���&����\��c*��:���
�����h��������\�^�E��e�e�e�e�g�f�W���
����_F��1�����0��
�
�'�+����&����	F��s1��2���_�u�u�<�9�1����,����_��~1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�g���������V��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�G���
����W'��^�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�;�4�1����Hù��l��h�����o������}���Y����R
��h^�����9�1��d��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��D�����
�d�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����0��
�d�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�I����P��S/��Dۊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�e��.����8����l��A�����u�u��
���W��^����F�D�����
�
�;�6�;�9�>��&����Z�=��*����
����u�BϺ�����O��N�����4�u�
�
�9�>����0����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��E���&�4�0���o��������l��T��!�����n�u�w�.����Y����f��V��4���g�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����,����_��~1�*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�֓�]��[��<��
�'�2�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��L�U���&�2�4�u����������lW��V�����;�&�2�o���;���:���F��P ��U���
�;�6�9�3��F܁�	����l��PN�&������o�w�m�L���Yӕ��]��G1�� ���4�0��
�c�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y����� �&�4�0���C�������`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�w�]�}�W�������lV��Y������d�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G���
����W'��Z�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��3��������9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������r/��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�e� �&�6�8�6���L����E
��^ �����u��
���f�W���
����_F��1�����0��
�`�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l*��^�����0�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h"�����;�7�0�
�%�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�M���I����V��^�E��n�u�u�&�0�<�W���&����G��V�����
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�>�4��������R��[
�����o������M���I��ƹF��^	��ʥ�`��2��:�)�G���&����	F��s1��2������u�f�}�������9F������%�`��2��0����	����	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�u�W�W���������h&�����<�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�B�������Z��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�>�5����&¹��l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��4��������C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��@���2��8�!�f�<�(���&����Z�=��*����n�u�u�$�:����&ƹ��T��Z��D���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�h�?���5����lT��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�B�������Z��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�<�=�>�4�(݁�	����l��D��Oʆ�����]�}�W�������lS��^	�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&������C1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ƹ��T��Z��F���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�`��:�;����Փ�C9��S1��*���u�u��
���L���Yӕ��]��G1��=����8�!�f�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l.��_"�����
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lS��^	�����
�
�'�2�m��3���>����v%��eN��@ʱ�"�!�u�|�m�}�G��I����V��^�N���u�&�2�4�w��(�������G9��V�����;�&�2�o���;���:���F��P ��U���
�<�=�<�>��(�������A��N��1�����o�u�g�f�W���
����_F��1�����8�!�`�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��=����8�!�`�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�L����[*��^��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�`��0�����L����E
��G��U����
���w�`�P���s���@��V��*ߊ�<�=�<�<����������g"��x)��*�����}�`�3�*����P���F��P ��U���
�<�=�<�>��(�������g"��x)��*�����}�`�3�*����P���V��^�E��e�e�e�n�w�}�����Ƽ�9��P�����c�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u����������9��h��*���2�o�����4��Y���9F������%�`��2��0��������TF��d:��9�������w�l�W������]ǻN�����9�%�`��0�����N����TF��d:��9�������w�l�W������F��L�E��e�e�e�e�g��}���Y����R
��h[�����<�<�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1����1����Z��hY�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��4��������Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u����������9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������2��8�#�e��������l��T��!�����n�u�w�.����Y����{��{�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�B�������Z��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����1����Z��hW�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�<�?�4����&����_��Y1���������W�W���������h&�����<�
�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&ƹ��T��Z��Dڊ�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��l.��_"�����e�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�h�?���5����lW��V�����;�&�2�o���;���:���F��P ��U���
�<�=�<�>��G���&����C��T��!�����u�h�p�z�}���Y����R
��h[�����<�<�
�d�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��@���2��8�!�f�����Cӵ��l*��~-��0����}�`�1� �)�W���C���V��^�E��e�e�n�u�w�.����Y����{��{����
�%�#�1�>�����Y����)��tUךU���<�;�9�%�b���������9��h��*���2�o�����4��Y���9F������%�`��2��0���&����Z�=��*����
����u�BϺ�����O��N�����4�u�
�
�>�5����&�ԓ�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*���=�<�<�
�e�<�(���&����Z�=��*����n�u�u�$�:����&ƹ��T��Z��D؊�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(�������G9��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����1����Z��h_�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�`��0�����H����l��h�����o������}���Y����R
��h[�����<�<�
�f�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l.��_"�����a�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9����9���!�d�
�'�0�g�$���5����l0��c!��]���1�"�!�u�~�g�W��I����V��^�E��u�u�&�2�6�}�(ځ�����^��Z�����1�<�
�<�w�}�#���6����9F������%�`��2��0���&����_��E��Oʆ�����m�}�G��Y����Z��[N��@���2��8�!�f���������g"��x)��*�����}�`�3�*����P���F��P ��U���
�<�=�<�>��B�������`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�w�]�}�W�������lS��^	�����
�`�4�
�;���������g"��x)��N���u�&�2�4�w��(�������G9��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�8�����I����@��N��1��������}�F�������V�=N��U���;�9�%�b��*����&ù��V�=��*����
����u�BϺ�����O�
N��E��e�e�e�e�g�m�L���Yӕ��]��G1��9���<�<�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1����5����^��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�b��*����&¹��l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��2�;����ד�A��N��1��������}�F�������V�S��E��e�e�e�e�g�m�U�ԜY�ƿ�T����*����8�!�d�6���������\��c*��:���n�u�u�&�0�<�W���&����Z��h_�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��2�;����ԓ�]9��PN�&���������W��Y����G	�UךU���<�;�9�%�`�� �������C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��B���"�<�<�
��-��������TF��d:��9����_�u�u�>�3�Ϯ�N������C1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�`�� �������Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u����������l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G���s���@��V��*݊�:��8�!�d�<�(���&����Z�=��*����n�u�u�$�:����&Ĺ��D*��^��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u����������l��D��Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�j�;�������9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"�<�<����������@��N��1�����_�u�w�4����	�ѓ�\��Z��A���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�j�;�������9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(���5����lS��E��Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��[���F��P ��U���
�:��8�#�h��������l��T��!�����n�u�w�.����Y����	��^��*ߊ�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(���5����lP��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�@�������G9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�b��"�<�>��(�������]9��PN�&������_�w�}����Ӗ��l*��{�����4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�@�������G9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(؁�����Z��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����F�D�����
�
�:��:�)�@���&����Z��^	��U���
���n�w�}�����Ƽ�9��@"�����
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(؁�����Z��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����5����^��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b��"�>�4�(ׁ�	����l��D��Oʆ�����]�}�W�������lQ��X�����m�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����5����^��1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&����Z��hW�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����l�N�����u�
�
�:��0��������W9��h��U����
���l�}�Wϭ�����C9��{�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����Z��h_�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&Ĺ��D*��^��E���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b��*����&�֓�C9��S1��*���u�u��
���L���Yӕ��]��G1��9���<�<�
�e�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l*��{����
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lQ��X�����d�
�'�2�m��3���>����v%��eN��@ʱ�"�!�u�|�m�}�G��I����V��^�N���u�&�2�4�w��(���5����lW��V�����;�&�2�o���;���:���F��P ��U���
�:��8�#�l�(�������A��N��1�����o�u�g�f�W���
����_F�� 1�����<�
�g�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��9���<�<�
�g�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�N������C1�*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�b�� �4����K����E
��G��U����
���w�`�P���s���@��V��*݊�:��8�!�f���������g"��x)��*�����}�`�3�*����P���F��P ��U���
�:��8�#�l�(�������g"��x)��*�����}�`�3�*����P���V��^�E��e�e�e�n�w�}�����Ƽ�9��@"�����f�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���������� 9��h��*���2�o�����4��Y���9F������%�b��"�>�4�(�������TF��d:��9�������w�l�W������]ǻN�����9�%�b�� �4����M����TF��d:��9�������w�l�W������F��L�E��e�e�e�e�g��}���Y����R
��hY�����8�!�d�
�'�+����&����	F��s1��2���_�u�u�<�9�1����5����^��Z�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��2�;�������Z��^	��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u����������9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y������"�<�<��h��������l��T��!�����n�u�w�.����Y����	��^��*���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�N���
����W*��^�����
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������l_��Y�����<�<��2������Cӵ��l*��~-��0����}�`�1� �)�W���C���V��^�E��e�e�n�u�w�.����Y����f��V��9���!�<�=�;�6���������\��c*��:���n�u�u�&�0�<�W���&����R
��{�����=�;�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�H¹��@��R
�����:��
�;�$�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��h_�� ���4�0��8�#�2�>������5��h"��<������}�b�9� ���Y���F�^�E��e�e�e�e�l�}�Wϭ�����C9��h;�����1�<�<�� �3��������l��T��!�����n�u�w�.����Y����l3��T�����<��"�;�6��������5��h"��<���h�r�r�_�w�}����Ӗ��9��R�����
�;�&�2�m��3���>����F�D�����
�g��0�%�4�������5��h"��<���h�r�r�_�w�}����Ӗ��9��R�����
�%�#�1�>�����Y����)��tUךU���<�;�9�%�f�����5����l��A�����u�u��
���W��^����F�D�����:�9������������lV�=��*����
����u�W������F��L�N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���&����r��B��F���3�
�f�
�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��U��4��� �
�f�e�%�:�E��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����:�9�'��#�h�(ށ�����Q�=��*����
����u�W������]ǻN�����9�4�'�7�8�����&�Փ�l��h\�G��������4���Y����\��XN�N���u�&�2�4�w�/�(�������F��1�����g�b�u�u���8���&����|4�N�����u�|�_�u�w�4��������\	��E�����
�
�0�
�f�o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1�����'� �
�f�b�/���A����`2��{!��6�����u�e�3�*����P���F��P ��U���
�:�9�'��)�B܁�&����W��T��!�����
����_�������V�=N��U���;�9�4�'�5�2�6�������lQ��R	��D��o������!���6�����Y��E��u�u�&�2�6�}��������A)��h[��M���2�g�e�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��[/��:���`�
�
�0��o�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V������'� �
�d�l�(���&����\��c*��:���
�����}�������9F������4�'�7�:��/����J����A��\�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�/����8����G9��h_�����g�g�u�u���8���&����|4�N�����u�|�_�u�w�4��������\	��E�����
�f�'�2�e�o�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����'��!�`��i����K����	F��s1��2������u�g�9� ���Y����F�D�����'�
�:�9�%����&�ӓ�V��]�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%���������lS��1��*��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������\	��E�����
�
�0�
�e�o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1�����'� �
�d�f�/���M����`2��{!��6�����u�e�3�*����P���F��P ��U���
�:�9�'��)�Bށ�&����T��T��!�����
����_�������V�=N��U���;�9�4�'�5�2�6�������lU��R	��G��o������!���6�����Y��E��u�u�&�2�6�}��������A)��h[��A���2�g�c�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��[/��:���`�
�
�0��o�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V������'� �
�f�k����K����	F��s1��2������u�g�9� ���Y����F�D�����'�
�:�9�%����&Ĺ��T9�� Y��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�?��������W��h��*��g�o�����4���:����V��X����n�u�u�&�0�<�W���&����r��B��D���'�2�g�m�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��X�����!�`�
�e�%�:�E��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����:�9�'��#�h�(�������_��N��1��������}�GϺ�����O��N�����4�u�'�
�8�1��������T��R	��F��o������!���6�����Y��E��u�u�&�2�6�}��������A)��h[��Dي�0�
�f�b�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��X�����
�d�d�
�2��D��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����:��'� ��l�Fځ�����Q�=��*����
����u�W������]ǻN�����9�4�'�7�8�����&�ߓ�l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}��������A)��hZ��E���2�g�g�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l��[/��:���a�
�
�0��n�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V������'� �
�n�o����K����	F��s1��2������u�g�9� ���Y����F�D�����'�
�:�9�%����&����T9��Y��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�?��������_��h��*��g�o�����4���:����V��X����n�u�u�&�0�<�W���&����r��B��L���'�2�g�a�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��X�����!�a�
�
�2��D��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����:��'� ��d�@�������F��d:��9�������w�m��������l�N�����u�'�
�:�;�/�8���Mʹ��A��]�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�/����8����G9��hW�����f�b�o����0���/����aF�
�����e�n�u�u�$�:��������\
��E!��*���d�
�0�
�d�o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1�����'� �
�l�f�����J���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�7�:��%�(�(���H����T9��\��U���
���
��	�%���Y����G	�UךU���<�;�9�4�%�?��������_��1����m�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����_'��x��Aӊ�a�'�2�g�n�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h������!�a�
�b�/���@����`2��{!��6�����u�e�3�*����P���F��P ��U���9�
�:�
�8�-�Fށ�����9��T��!�����
����_�������V�=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����c�o�����}���Y����R
��{1��*���
�:�%�&�%�:�A��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����;�b�3�
�d�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������:�
�:�%�f���������l��T��!�����
����_������\F��d��Uʦ�2�4�u�8��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʼ�
�!��'��2�(���	����F9��1��G��������4���Y����W	��C��\�ߊu�u�<�;�;�4�(���?����\	��^����� �b�l�%�e�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������[1��*���
�:�%�g��5�(���A�Г� T�=��*����
����u�W������]ǻN�����9�7�:�
�#���������l��h��M���%�g�o����0���/����aF�
�����e�n�u�u�$�:��������G9��E1�����c�%�<�3��d�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*����0�'�<�>���������U��V��G��������4���Y����\��XN�N���u�&�2�4�w�/�(���?����\	��Y��@���
�f�u�u���8���&����|4�N�����u�|�_�u�w�4��������G9��E1�����b�e�3�
�d�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*����'��:��j�Fځ�&���� R�=��*����
����u�W������]ǻN�����9�4�'�9��2�(���	����S��h��G��o������!���6�����Y��E��u�u�&�2�6�}��������l*��G1�*���f�3�
�a�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��C1�����:�
�b�d�����O����g"��x)��*�����}�u�8�3���B�����Y�����9�
�:�
�8�-�E؁�L�ӓ�F9��N�&���������W������\F��d��Uʦ�2�4�u�'��)�1���5����Q��1�����`�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�����u	��{��*���d�
�
� �e�e�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�g��h�O���&����	F��s1��2������u�g�9� ���Y����F�D�����'�
�!��%�����N����
9��h\�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�/��������\�� 1�*���3�
�b�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l
��q��9���
�b�d�
�f�;�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����!��'��8��@��&�ԓ�F9��N�&���������W������\F��d��Uʦ�2�4�u�'��)�1���5����Q��1�*���g�g�o����0���/����aF�
�����e�n�u�u�$�:��������l ��h"����
�`�d�
�"�o�A��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��B��&����
V�=��*����
����u�W������]ǻN�����9�4�'�9��2�(���	����S��B1�A��������4���Y����\��XN�N���u�&�2�4�w�/�(���?����\	��W��*���d�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�g�
�`�f�;�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����!��'��8��N��&����lU��T��!�����
����_�������V�=N��U���;�9�4�'�;���������
9��h]�� ��c�o�����4���:����V��X����n�u�u�&�0�<�W���&����\��X��Gӊ�`�a�3�
�f�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��3����:�
�l�f��(���J���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�9�
�:��2���&�ӓ�l ��_�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%���������C9��h_��B���
�g�u�u���8���&����|4�N�����u�|�_�u�w�4��������G9��E1�����l�d�
�
�"�n�A��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e��B�������F��d:��9�������w�m��������l�N�����u�'�
�!��/�;���&�ߓ�9��h��F��o������!���6�����Y��E��u�u�&�2�6�}��������l*��G1�*���d�
� �f�o�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��[�����:�%�g�
�b�l�(���J���5��h"��<������}�w�2����I��ƹF��^	��ʴ�'�9�
�:��2���&�ӓ� 9��h]�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�/��������\��1�*���3�
�`�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��l
��q��9���
�l�d�
�b�;�(��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*��� �!�`�&�1��A���	���5��h"��<������}�b�9� ���Y����F�D�����
�0� �!�a�.����O�֓�Q�=��*����
����u�BϺ�����O��N�����4�u�:�9�/�	�8���OĹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�2�(��� ����Q��C�����e�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӄ��_9��c����
� �d�c��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h=��0��� �
�l�3��m�F���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����7�:��'�"��N�������U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}��������F��1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������K*��x��A܊� �d�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q	��h �����'�
�a�3��n�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����;�1�
�0�:�n�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�&�1��@���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʴ�
��3�8�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�l��h��*��e�o�����}���Y����R
��G1�����1�d�b�u�w��;���B�����Y�����<�
�1�
�f�}�W���5����9F������4�
�<�
�3��@��;����r(��N�����4�u�%�&�0�?���M����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:����	����l��h_�U������n�w�}�����ƭ�l��h��*���u�u����f�W���
����_F��h��*���
�c�u�u���6��Y����Z��[N��*���
�1�
�b�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��k�MϜ�6����l�N�����u�%�&�2�5�9�B���Y����v'��=N��U���;�9�4�
�>�����M����|)��v �U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�<�(���&����T�,��9���n�u�u�&�0�<�W���
����W��N�7�����_�u�w�4��������T9��S1�E������]�}�W�������C9��P1����l�o�����}���Y����R
��G1�����1�d�m�o���2���s���@��V�����2�7�1�a�f�g�5���<����F�D�����%�&�2�7�3�h�G��;����r(��N�����4�u�%�&�0�?���H����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lT��T��:����n�u�u�$�:����	����l��h\�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�e�u�u���6��Y����Z��[N��*���
�1�
�d�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����W��N��:����_�u�u�>�3�Ͽ�&����Q��\�Oʗ����_�w�}����Ӈ��@��U
��G���o�����W�W���������D�����g�a�o����9�ԜY�ƿ�T�������7�1�g�f�m��8���7���F��P ��U���&�2�7�1�e�o�MϜ�6����l�N�����u�%�&�2�5�9�E��CӤ��#��d��Uʦ�2�4�u�%�$�:����J���$��{+��N���u�&�2�4�w�-��������R�,��9���n�u�u�&�0�<�W���
����W��]��U�����n�u�w�.����Y����Z��S
��A���u����l�}�Wϭ�����R��^	�����`�u�u����L���Yӕ��]��V�����1�
�c�u�w��;���B�����Y�����<�
�1�
�a�}�W���5����9F������4�
�<�
�3��C���Y����v'��=N��U���;�9�4�
�>�����L����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�L������]�}�W�������C9��P1����m�o�����}���Y����R
��G1�����1�f�b�o���2���s���@��V�����2�7�1�a�a�g�5���<����F�D�����%�&�2�7�3�i�B��;����r(��N�����4�u�%�&�0�?���I����|)��v ���2�;�_�_�w�}�Z����Ư�A��CN�����}�%��
�$�t�����ƿ�R��Z�����u�x�u�u�6��$�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���6���&�u�h�4��	��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����YNךU���u�u�u�u�w�}�W���	����U��S�����
�&�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���&�4�0�����������TF��D��U���6�&�{�x�]�}�W���&����R
��v'��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����f��V��4���
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^�����<�
�1�
�b�t����Y���F�N��U���u�u�u�u�w��(�������r/��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�u�w�}�W�������C9��P1����|�!�0�u�w�}�W���Y���F�N��U���
�
�;�6�;�9�>�������W9��R	��Hʥ�e� �&�4�2��(߁�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g���������9��R	�����;�%�:�0�$�}�Z���YӖ��l3��T�����e�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��@��R
��*ڊ�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϮ�I����P��S/��E���
�9�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\���!�0�u�u�w�}�W���Y���F���*���6�9�1��g�-����DӖ��l3��T�����e�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h^�����9�1��d��-����	����R��P �����&�{�x�_�w�}�(߁�����V��h_�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�]��[��<��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^�����<�
�1�
�b�t����Y���F�N��U���u�u�u�u�w��(�������r/��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����g�|�!�0�w�}�W���Y���F�N��U���u�
�
�;�4�1����Hù��l��h����u�
�
�;�4�1����Hù��l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�G���
����W'��^�����4�&�2�u�%�>���T���F��1�����0��
�e�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��b ������
�e�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R
��v'��E���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�;�4�1����Hù��V�
N��E���&�4�0���m�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�;�4�1����H¹��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��b ������
�d�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���6�9�1��f���������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��D�����
�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�����V��h_�����9�
�'�2�k�}�(߁�����V��h_�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��Y������d�
�'�0�<����Y����V��C�U���%�e� �&�6�8�6���H����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�e� �&�4�2��(���	����[��G1�����9�d�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����0��
�d�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(߁�����V��h_�����u�h�%�e��.����8����l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����V��h_�����9�
�'�2�6�.��������@H�d��Uʥ�e� �&�4�2��(�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�9�>����0����R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}��������T9��S1�A���=�;�_�u�w�}�W���Y���F�N����� �&�4�0���E���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9��b ������
�g�4��1�(������C9��b ������
�g�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�;�6�9�3��F݁�����@��YN�����&�u�x�u�w�-�G���
����W'��\�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�m�"�������z9��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e� �&�6�8�6���K����E
��G�����_�u�u�u�w�}�W���Y���C9��b ������
�g�%�2�}�JϮ�I����P��S/��D��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��b ������
�f�4��1�(���Ӈ��Z��G�����u�x�u�u�'�m�"�������z9��h�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����R
��v'��F���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y����������7�1�l�a�w�5��ԜY���F�N��U���u�u�u�%�g���������U��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��Uʥ�e� �&�4�2��(�������W9��R	��Hʥ�e� �&�4�2��(�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������lW��G��U���<�;�%�:�2�.�W��Y����lV��Y������d�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l3��T�����d�
�'�2�k�}��������EW��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�G���
����W'��]�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e� �&�4�2��(���	����[��h^�����9�1��d�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(�������W9��R	�����;�%�:�0�$�}�Z���YӖ��l3��T�����d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����0��
�a�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�%�&�0�?���M�Ƹ�V�N��U���u�u�u�u�w�}�W���	�֓�]��[��<��
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�d�d�}����s���F�N��U���u�u�u�u�'�m�"�������z9��h�����%�0�u�h�'�m�"�������z9��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����f��V��4���a�%�0�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��Fہ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�;�6�9�1��l�(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��Y������d�
�%�!�9�^������F�N��U���u�u�u�u�'�m�"�������z9��h����u�
�
�;�4�1����H��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�"�������z9��h�����%�0�u�&�>�3�������KǻN��*ڊ�;�6�9�1��l�(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e� �&�6�8�6���L����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_���
����W��Z�����u�u�u�u�w�}�W���Y���F���*���6�9�1��f���������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����H���G��d��U���u�u�u�u�w�}�W���YӖ��l3��T�����d�
�%�#�3�-����DӖ��l3��T�����d�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���&�4�0���h����Y����T��E�����x�_�u�u����������lW��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��3��������9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�;�6�9�3��Fځ�	����O�C��U���u�u�u�u�w�}�W���YӖ��l3��T�����d�
�'�2�k�}�(߁�����V��h_����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l3��T�����d�4�
�9��/�Ͽ�
����C��R��U���u�u�%�e��.����8����R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�m�"�������z9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������C9��P1����a�u�=�;�]�}�W���Y���F�N��U���%�e� �&�6�8�6���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR�����ߊu�u�u�u�w�}�W���Y���F��1�����0��
�
�'�+���������h;�����1��d�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�;�6�9�3��F����ƭ�@�������{�x�_�u�w��(�������r/��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g���������9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�;�6�9�3��F���&����O��_�����u�u�u�u�w�}�W���Y����f��V��4���
�'�2�i�w��(�������r/��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*؊�%�#�1�%�2�}����Ӗ��P��N����u�
�
�;�4�1����K����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��3��������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���Y���F�N��U���
�;�6�9�3��E���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lV��Y������g�4�
�;�����E�Ƽ�9��D�����
�
�%�#�3�W�W���Y���F�N��Uʰ�1�<�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���&�4�0�����������]F��X�����x�u�u�%�g���������9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�9�>����0�ԓ�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��E���&�4�0����������G��d��U���u�u�u�u�w�}�WϮ�I����P��S/��G���0�u�h�%�g���������]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����,����_��~1�����9�
�'�2�6�.��������@H�d��Uʥ�e� �&�4�2��(܁�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�e� �$�<����&����l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�Wǿ�&����Q��[�U���;�_�u�u�w�}�W���Y���F�N��E���&�4�0�����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����O����[��=N��U���u�u�u�u�w�}�W���Y����f��V��4���
�%�#�1�'�8�W��	�֓�]��[��<���4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h^�����9�1��f�'�8�W�������A	��D�X�ߊu�u�
�
�9�>����0�Փ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e� �&�6�8�6���&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h^�����9�1��f�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(߁�����V��h]�����i�u�
�
�9�>����0����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������r/��h�����%�0�u�&�>�3�������KǻN��*ڊ�;�6�9�1��i��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�;�6�;�9�>�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������l_��N�����u�u�u�u�w�}�W���Y���F��h^�����9�1��a�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��Y����l�N��U���u�u�u�u�w�}�WϮ�I����P��S/��A���
�9�
�'�0�a�W���&����R
��v'��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��b ������
�
�'�0�<����Y����V��C�U���%�e� �&�6�8�6���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�;�6�9�3��C��������T�����d�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��b ������
�
�%�!�9�^������F�N��U���u�u�u�u�'�m�"�������z9��G��U��%�e� �&�6�8�6���B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�g���������9��h��*���2�4�&�2�w�/����W���F�G1�� ���4�0��
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N����� �&�4�0���(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9��b ������
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�e�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�����V��h[�����1�%�0�u�j�-�G���
����W'��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l3��T�����`�%�0�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��B�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��E���&�4�0�������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l3��T�����`�4�
�9�~�t����Y���F�N��U���u�u�u�
��3��������l��PN�U���
�;�6�9�3��B�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�9�>����0�Г�C9��S1�����&�<�;�%�8�8����T�����h;�����1��c�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���6�9�1��a�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�%�$�:����@���G��d��U���u�u�u�u�w�}�W���YӖ��l3��T�����c�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�f�}����s���F�N��U���u�u�u�u�'�m�"�������z9��V�����'�2�i�u����������lP��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*܊�'�2�4�&�0�}����
���l�N��E���&�4�0�����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^�����9�1��c�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ù��@��R
��*܊�%�#�1�|�w�5��ԜY���F�N��U���u�%�e� �$�<����&Ź��V�
N��E���&�4�0���f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�e� �&�6�8�6���&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��D�����
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����0��
�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ù��@��R
��*݊�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�d�e�w�5��ԜY���F�N��U���u�u�u�%�g���������9��h��*���2�i�u�
��3��������l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��v'��*���2�4�&�2�w�/����W���F�G1�� ���4�0��
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h;�����1��b�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R
��v'��*���#�1�|�u�?�3�}���Y���F�N��U���%�e� �&�6�8�6���&����Z�G1�� ���4�0��
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e� �&�4�2��(ׁ�	����l��PN�����u�'�6�&�y�p�}���Y����f��V��4���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��b ������
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����4�
�<�
�3��B�������9F�N��U���u�u�u�u�w�}�W���&����R
��v'��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����UF��G1�����1�d�l�u�?�3�}���Y���F�N��U���u�u�%�e��.����8����R��[
�����i�u�
�
�9�>����0�ޓ�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����V��hV�����4�&�2�u�%�>���T���F��1�����0��
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��Y������m�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(߁�����V��hV�����1�|�u�=�9�W�W���Y���F�N��Uʥ�e� �&�4�2��(ׁ����F��1�����0��
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C���� �&�4�0���(�������A��V�����'�6�&�{�z�W�W���&ù��@��R
��*ӊ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��D�����
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�����V��hW�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����d�m�u�=�9�W�W���Y���F�N��U���u�%�e� �$�<����&ʹ��l��h����u�
�
�;�4�1����@����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(�������r/��h��ʴ�&�2�u�'�4�.�Y��s���C9��b ������
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l3��T�����l�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������r/��h�����|�u�=�;�]�}�W���Y���F�N����� �&�4�0���(������C9��b ������
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��Dۊ�;�6�9�1�>�4�;�������E
��G��U���<�;�%�:�2�.�W��Y����lW��b ������8�!�:����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�d�
�;�6�;�9����5����l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���Y���F�N��U���d� �&�4�2���������R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hZ�\ʡ�0�u�u�u�w�}�W���Y���F�N��*��� �&�4�0��0����0����l��h����u�
�d� �$�<��������D/��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	����f��V��9���!�:��
�%�:�����Ƽ�\��D@��X���u�%�d�
�9�>��������\��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�f���������^��X��*���2�i�u�%�4�3����HŹ��9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�d��3��������G*��~ �����1�|�u�=�9�W�W���Y���F�N��Uʥ�d�
�;�6�;�9����5����l��PN�U���d� �&�4�2���������9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�F݁�����Z��h�����%�0�u�&�>�3�������KǻN��*����0�'�<�>���������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�d�
�9�4��0����&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��-��������R�C��U���u�u�u�u�w�}�W���Y�����1�����<�<�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�h�G������F�N��U���u�u�u�u�w�}���&����A*��^�����1�%�0�u�j�-�F݁�����Z��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����l%��V�����%�0�u�&�>�3�������KǻN��*����0�'�<�>���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h_��6���'�<�<�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&�ԓ�_��{�����
�9�|�|�#�8�W���Y���F�N��U���u�
�g��2�/����&����Z�G1�*���4��8�!�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�<�<�<�9�?����	����l��PN�����u�'�6�&�y�p�}���Y������C�����1�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h"�����;�7�0�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&¹��^��r �����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�m�~�)����Y���F�N��U���u�u�u�u����������_��V�����'�2�i�u����������_��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ד�Z��^+�����
�'�2�4�$�:�W�������K��N������8�!��6�1��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��D���8�!��4�;�9����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��Z��0���9�1�4�
�;�t�^Ϫ���ƹF�N��U���u�u�u�u����������_��G��U��%�d��8�#��������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������9��h��*���2�4�&�2�w�/����W���F�G1��=����8�!�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�<�=�<�<����������TF������!�9�2�6�g�W�W���Y���F��DךU���u�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��P�����e�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�n�t����Y���F�N��U���u�u�u�u�w��(�������G9��V�����'�2�i�u����������9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����[*��^��*���2�4�&�2�w�/����W���F�G1��=����8�!�e�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9����9���!�e�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�����^��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�<�=�<�>��(������C9����9���!�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���=�<�<�
�g�<�(���&������^	�����0�&�u�x�w�}����1����Z��h_�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ӓ�Z��^��*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�l�c�}����s���F�N��U���u�u�u�u�'�h�?���5����lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�<�=�>�4�(�������W9��R	��Hʥ�`��2��:�)�F߁�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�b���������9��R	�����;�%�:�0�$�}�Z���YӖ��l.��_"�����e�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ƹ��T��Z��Dڊ�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�b���������9��h��\���!�0�u�u�w�}�W���Y���F���*���=�<�<�
�g�-����DӖ��l.��_"�����e�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h[�����<�<�
�d�6���������@��YN�����&�u�x�u�w�-�B�������Z��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�L����[*��^��D���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y����������7�1�l�a�w�5��ԜY���F�N��U���u�u�u�%�b���������9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��M���!�0�u�u�w�}�W���Y���F�N��U���
�<�=�<�>��F���&����C��R������2��8�#�l�(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�`��:�;�������C�������%�:�0�&�w�p�W���	�ӓ�Z��^��*���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&������C1�*���2�i�u�%�4�3����HŹ��9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�`��:�;�������R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h[�����<�<�
�d�'�8�W��	�ӓ�Z��^��*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h&�����<�
�g�4��1�(���Ӈ��Z��G�����u�x�u�u�'�h�?���5����lW��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����1����Z��h_�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF��G1�����1�l�a�u�?�3�}���Y���F�N��U���u�u�%�`��:�;�������R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ߊ�<�=�<�<��o��������V�
N��@���2��8�!�f��������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`��0�����H����V��D��ʥ�:�0�&�u�z�}�WϮ�L����[*��^��G���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�����^��\�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`��0�����H����l��G�����u�u�u�u�w�}�W���Y�����h&�����<�
�g�%�2�}�JϮ�L����[*��^��G�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lS��^	�����
�f�4�
�;���������]F��X�����x�u�u�%�b��������� 9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�B�������Z��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����l�a�u�=�9�W�W���Y���F�N��U���u�%�`��0�����H����l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��Y�����u�u�u�u�w�}�W���Y���F���*���=�<�<�
�d�<�(���&����Z�G1��=����8�!�d��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�`��2��0���&������^	�����0�&�u�x�w�}����1����Z��h_�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������G9��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`��2��0���&����_�N�����u�u�u�u�w�}�W���Y����lS��^	�����
�f�%�0�w�`����1����Z��h_����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l.��_"�����a�4�
�9��/�Ͽ�
����C��R��U���u�u�%�`��:�;�������R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�h�?���5����lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������C9��P1����a�u�=�;�]�}�W���Y���F�N��U���%�`��2��0���&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lU��N�����u�u�u�u�w�}�W���Y���F��h[�����<�<�
�a�6��������F��1�����8�!�d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�`��2��:�)�Fہ�����@��YN�����&�u�x�u�w�-�B�������Z��1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u����������R��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`��2��:�)�Fہ�	����O�C��U���u�u�u�u�w�}�W���YӖ��l.��_"�����a�%�0�u�j�-�B�������Z��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�Z��^��*���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�`��0�����Hƹ��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b���������9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Yۇ��@��U
��L��u�=�;�_�w�}�W���Y���F�N��Uʥ�`��2��:�)�Fځ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������S�C��U���u�u�u�u�w�}�W���Y�����h&�����<�
�`�4��1�(������C9����9���!�d�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����2��8�#�l�(���Ӈ��Z��G�����u�x�u�u�'�h�?���5����lW��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��4��������l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������2��8�#�l�(������F��R ��U���u�u�u�u�w�}�W���	�ӓ�Z��^��*���%�0�u�h�'�h�?���5����lW��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����[*��^��*���#�1�%�0�w�.����	����@�CךU���
�
�<�=�>�4�(ށ�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�`��0�����H����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_���
����W��Z�����u�u�u�u�w�}�W���Y���F���*���=�<�<�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���@�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ӓ�Z��^��*ۊ�%�#�1�%�2�}�JϮ�L����[*��^��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9����9���!�d�%�0�w�.����	����@�CךU���
�
�<�=�>�4�(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�<�=�<�<������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l.��_"�����
�%�#�1�~�}����s���F�N��U���u�u�%�`��:�;����ד�A��S��*ߊ�<�=�<�<��f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�`��2��0��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l.��_"�����
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9����9���!�g�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����%�&�2�7�3�d�C������F�N��U���u�u�u�u�w�}����1����Z��h\�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����g�m�u�=�9�W�W���Y���F�N��U���u�%�`��0�����K����E
��G��U��%�`��2��0��������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������9��R	�����;�%�:�0�$�}�Z���YӖ��l.��_"�����
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�L����[*��^��*���2�i�u�%�4�3����HŹ��9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�`��:�;����ԓ�C9��SG��U���;�_�u�u�w�}�W���Y���F��1�����8�!�g�%�2�}�JϮ�L����[*��^��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��P�����f�4�
�9��/�Ͽ�
����C��R��U���u�u�%�`��:�;����Փ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���������� 9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Yۇ��@��U
��L��u�=�;�_�w�}�W���Y���F�N��Uʥ�`��2��:�)�D���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9����9���!�f�4�
�;�����E�Ƽ�9��P�����f�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���=�<�<�
��/�Ͽ�
����C��R��U���u�u�%�`��:�;����Փ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�`��2��0����	����[��G1�����9�d�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����8�!�f�4��1�^�������9F�N��U���u�u�u�u�w��(�������G9��G��U��%�`��2��0���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��4��������R��[
�����4�&�2�u�%�>���T���F��1�����8�!�a�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���=�<�<�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����L����[��=N��U���u�u�u�u�w�}�W���Y����{��{�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�g�~�)����Y���F�N��U���u�u�u�u����������9��h��*���2�i�u�
��4��������R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����1����Z��hZ�����4�&�2�u�%�>���T���F��1�����8�!�a�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��P�����a�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������G9��V�����|�!�0�u�w�}�W���Y���F�N��*ߊ�<�=�<�<������E�Ƽ�9��P�����a�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h[�����<�<�
�
�'�+�����ƭ�@�������{�x�_�u�w��(�������G9��V�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����1����Z��h[�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��h��*���
�`�|�!�2�}�W���Y���F�N��U���u�u�
�
�>�5����&ƹ��l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��[�����u�u�u�u�w�}�W���Y���F���*���=�<�<�
��-����	����[��h[�����<�<�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�`��2��:�)�B����ƭ�@�������{�x�_�u�w��(�������G9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��4��������C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ߊ�<�=�<�<���������G��d��U���u�u�u�u�w�}�WϮ�L����[*��^��*���2�i�u�
��4��������9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�B�������Z��h�����%�0�u�&�>�3�������KǻN��*ߊ�<�=�<�<����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`��2��:�)�A���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��-��������R�C��U���u�u�u�u�w�}�W���Y�����h&�����<�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�o�C������F�N��U���u�u�u�u�w�}����1����Z��hX�����1�%�0�u�j�-�B�������Z��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����{��{�����%�0�u�&�>�3�������KǻN��*ߊ�<�=�<�<����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h[�����<�<�
�
�%�:�K���	����@��A_��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�L����[*��^��*���#�1�|�u�?�3�}���Y���F�N��U���%�`��2��0����	����[��h[�����<�<�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C�����2��8�#�j��������V��D��ʥ�:�0�&�u�z�}�WϮ�L����[*��^��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����{��{�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�l�c�}����s���F�N��U���u�u�u�u�'�h�?���5����lQ��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��G��u�=�;�_�w�}�W���Y���F�N��Uʥ�`��2��:�)�@���&����C��R������2��8�#�j������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�>�5����&Ĺ��V��D��ʥ�:�0�&�u�z�}�WϮ�L����[*��^��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�B�������Z��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�`��2��0��������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�9��P�����b�%�0�u�j�-�B�������Z��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ƹ��T��Z��M���
�9�
�'�0�<����Y����V��C�U���%�`��2��0��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�>�5����&˹��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�Wǿ�&����Q��[�U���;�_�u�u�w�}�W���Y���F�N��@���2��8�!�o�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����O����[��=N��U���u�u�u�u�w�}�W���Y����{��{�����4�
�9�
�%�:�K���&ƹ��T��Z��M���
�9�n�u�w�}�W���Y���F���U���_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h&�����<�
�
�'�0�<����Y����V��C�U���%�`��2��0����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������2��8�#�e����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��P�����m�4�
�9�~�t����Y���F�N��U���u�u�u�
��4��������C��R������2��8�#�e�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�<�?�4����&����_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��P�����l�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h&�����<�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����4�
�<�
�3��B�������9F�N��U���u�u�u�u�w�}�W���&������C1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�b�|�!�2�}�W���Y���F�N��U���u�u�
�
�>�5����&ʹ��l��h����u�
�
�<�?�4����&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h�?���5����l_��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��P�����l�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ƹ��T��Z��L���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��4��������R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h[�����<�<�
�
�%�:�K���&ƹ��T��Z��L�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��X�����e�4�
�9��/�Ͽ�
����C��R��U���u�u�%�b��*����&ù��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�� �������R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}��������T9��S1�A���=�;�_�u�w�}�W���Y���F�N������"�<�<����������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����J���G��d��U���u�u�u�u�w�}�W���YӖ��l*��{�����4�
�9�
�%�:�K���&Ĺ��D*��^��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��{�����
�
�'�2�6�.��������@H�d��Uʥ�b��"�<�>��(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*����8�!�e�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��D*��^��*���#�1�|�u�?�3�}���Y���F�N��U���%�b��"�>�4�(߁����F�� 1�����<�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��B���"�<�<�
�g�<�(���&������^	�����0�&�u�x�w�}����5����^��^�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��D*��^��E���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y����������7�1�l�a�w�5��ԜY���F�N��U���u�u�u�%�`�� �������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�A���=�;�_�u�w�}�W���Y���F�N������"�<�<��m��������V�
N��B���"�<�<�
�g�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�:��0���&������^	�����0�&�u�x�w�}����5����^��^�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�;�������V��E��I���%�6�;�!�;�l�(��Y���F�N�����u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�b��"�<�>��G���&����O��_�����u�u�u�u�w�}�W���Y����	��^��*���%�0�u�h�'�j�;�������V��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����Z��h_�����9�
�'�2�6�.��������@H�d��Uʥ�b��"�<�>��F���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�:��0���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��9���<�<�
�d�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��D*��^��D���
�9�
�'�0�a�W���&����Z��h_�����9�n�u�u�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lQ��X�����d�
�'�2�6�.��������@H�d��Uʥ�b��"�<�>��F�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���"�<�<�
�f�-����DӇ��P	��C1��D܊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����	��^��*���4�
�9�|�~�)����Y���F�N��U���u�u�
�
�8�����H¹��V�
N��B���"�<�<�
�f�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�:��:�)�F݁�	����l��PN�����u�'�6�&�y�p�}���Y����	��^��*���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��X�����d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�����Z��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����a�|�!�0�w�}�W���Y���F�N��U���u�
�
�:��0���&����_��E��I���
�
�:��:�)�F݁�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`�� �������l��PN�����u�'�6�&�y�p�}���Y����	��^��*���%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����Z��h_�����u�h�4�
�8�.�(���O����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�8�����H����l��G�����u�u�u�u�w�}�W���Y�����h"��9���!�d�
�'�0�a�W���&����Z��h_����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l*��{����
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
�8�����H����l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�`�� �������l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���Y���F�N��U���
�:��8�#�l�(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��X�����d�
�%�#�3�-����DӖ��l*��{����
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��9���<�<�
�f�'�8�W�������A	��D�X�ߊu�u�
�
�8�����H����V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�:��:�)�F܁����F��h�����#�c�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h"��9���!�d�
�%�!�9�^������F�N��U���u�u�u�u�'�j�;�������U��E��I���
�
�:��:�)�F��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��*����&�ғ�C9��S1�����&�<�;�%�8�8����T�����h"��9���!�d�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��9���<�<�
�a�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�%�&�0�?���M�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�\��Z��Dފ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�a�e�w�5��ԜY���F�N��U���u�u�u�%�`�� �������l��A�����u�h�%�b��*����&�ғ�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(؁�����Z��1�����&�<�;�%�8�8����T�����h"��9���!�d�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l*��{����
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�;�������R��G1�����u�=�;�_�w�}�W���Y���F�N��B���"�<�<�
�c�-����DӖ��l*��{����n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����<�
�`�4��1�(���Ӈ��Z��G�����u�x�u�u�'�j�;�������S��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�����Z��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����l�a�u�=�9�W�W���Y���F�N��U���u�%�b�� �4����L����E
��G��U��4�
�:�&��2����B���F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��9���<�<�
�`�6��������F�� 1�����<�
�`�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�:��8�#�l�(���Ӈ��Z��G�����u�x�u�u�'�j�;�������S��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b��*����&�ӓ�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���"�<�<�
�b�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����Z��h_�����u�h�%�b��*����&����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(���5����lW��G1�����0�u�&�<�9�-����
���9F���*����8�!�d�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�:��8�!�f�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�%�$�:����@���G��d��U���u�u�u�u�w�}�W���YӖ��l*��{�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�a�~�)����Y���F�N��U���u�u�u�u����������l��A�����u�h�%�b��*����&¹��l��d��U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@�������G9��G��U���<�;�%�:�2�.�W��Y����lQ��X�����d�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��D*��^��*���2�i�u�%�4�3����HŹ��9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�b��*����&¹��l��G�����u�u�u�u�w�}�W���Y�����h"��9���!�d�%�0�w�`����5����^��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ѓ�\��Z��G���
�9�
�'�0�<����Y����V��C�U���%�b��"�>�4�(݁�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�b�� �4����&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��9���<�<�
�
�'�+���������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�D��Y����l�N��U���u�u�u�u�w�}�WϮ�N������C1�����9�
�'�2�k�}�(؁�����Z��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����	��^��*؊�'�2�4�&�0�}����
���l�N��B���"�<�<�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h"��9���!�g�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�����Z��h�����|�u�=�;�]�}�W���Y���F�N������"�<�<������E�Ƽ�9��@"�����n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�����<�
�
�%�!�9����Y����T��E�����x�_�u�u����������l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���5����lU��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*���|�!�0�u�w�}�W���Y���F�N��U���
�
�:��:�)�D���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������O��_�����u�u�u�u�w�}�W���Y���C9��{�����
�
�%�#�3�-����DӖ��l*��{�����4�
�9�n�w�}�W���Y���F�N�����3�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hY�����8�!�f�%�2�}����Ӗ��P��N����u�
�
�:��0����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������"�<�<������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��l*��{�����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�8�����J����TF���*����8�!�f�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�:��8�#�i��������V��D��ʥ�:�0�&�u�z�}�WϮ�N������C1�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�\��Z��A���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y����������7�1�l�a�w�5��ԜY���F�N��U���u�u�u�%�`�� �������R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h]�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�:��8�!�c�<�(���&����Z�G1��9���<�<�
�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b��"�<�>��(���Ӈ��Z��G�����u�x�u�u�'�j�;�������9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�8�����M����TF������!�9�d�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��9���<�<�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�@�������G9��G��U��%�b��"�>�4�(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b��*����&ƹ��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��{�����
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1�����<�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����4�
�<�
�3��B�������9F�N��U���u�u�u�u�w�}�W���&����Z��h[�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����f�l�u�=�9�W�W���Y���F�N��U���u�%�b�� �4����&����_��E��I���
�
�:��:�)�B���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��2�;����ӓ�A��V�����'�6�&�{�z�W�W���&Ĺ��D*��^��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�@�������G9��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�:��:�)�B���&����O��_�����u�u�u�u�w�}�W���Y����	��^��*ߊ�'�2�i�u����������l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(؁�����Z��h�����%�0�u�&�>�3�������KǻN��*݊�:��8�!�a�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�:��8�#�k��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��X�����c�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�o�t����Y���F�N��U���u�u�u�u�w��(���5����lP��G1�����0�u�h�%�`�� �������R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����5����^��1�����&�<�;�%�8�8����T�����h"��9���!�c�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����	��^��*܊�'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�`�� �������R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��hY�����8�!�c�%�2�}�JϮ�N������C1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l*��{�����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�b�� �4����&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b��*����&Ĺ��l��h����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�4�Wǿ�&����Q��[�U���;�_�u�u�w�}�W���Y���F�N��B���"�<�<�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���N�Ƹ�V�N��U���u�u�u�u�w�}�W���	�ѓ�\��Z��B���
�9�
�'�0�a�W���&����Z��hY�����1�_�u�u�w�}�W���Y���F��SN��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��@"�����
�'�2�4�$�:�W�������K��N������"�<�<����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hY�����8�!�b�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����Z��hY�����1�|�u�=�9�W�W���Y���F�N��Uʥ�b��"�<�>��(������C9��{�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��9���<�<�
�
�'�+�����ƭ�@�������{�x�_�u�w��(���5����l^��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�����Z��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y���R��^	�����`�|�!�0�w�}�W���Y���F�N��U���u�
�
�:��0��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����V�����ߊu�u�u�u�w�}�W���Y���F�� 1�����<�
�
�%�!�9����Y����lQ��X�����m�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*����8�!�m�'�8�W�������A	��D�X�ߊu�u�
�
�8�����A����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b��"�<�>��(������R��X ��*���c�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lQ��X�����m�4�
�9�~�t����Y���F�N��U���u�u�u�
��2�;����ޓ�A��S��*݊�:��8�!�o�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�:��:�)�N���&����C�������%�:�0�&�w�p�W���	�ѓ�\��Z��L���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l*��{�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�l�c�}����s���F�N��U���u�u�u�u�'�j�;�������
9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��D���!�0�u�u�w�}�W���Y���F�N��U���
�:��8�#�d��������V�
N��B���"�<�<�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b��"�>�4�(ց�����@��YN�����&�u�x�u�w�-�@�������G9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��2�;����ߓ�A��S�����;�!�9�d��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B���"�<�<�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����5����^��1�����h�%�b�� �4����B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�n���������Z��P��*���#�1�%�0�w�.����	����@�CךU���
�
�;�6�;�9����1����]9��h��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�N���
����W*��^�����
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^�����<�
�1�
�b�t����Y���F�N��U���u�u�u�u�w��(���������C&�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�m�~�)����Y���F�N��U���u�u�u�u����������^��^	�����
�9�
�'�0�a�W���&����R
��{�����=�;�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ӊ�;�6�9�1�>�4�?���0����V��D��ʥ�:�0�&�u�z�}�WϮ�@����P��S"�����2��
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l3��T�����<��2���/���Y����\��h��C��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ�]��[������2��
�'�+����Y����l�N��U���u�u�u�u�w�-�N���
����W*��^�����
�'�2�i�w��(���������C&�����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����[�����:�%�&�'�0�k�FϿ�
����C��R��U���u�u�<�
�>���������A��W�����2�
�'�6�m�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Yӏ����D�����d�b�|�!�2�}�W���Y���F�N��U����9�
�:��2��������
W�
N��*����'��:��l����J�ד�]ǻN��U���u�u�u�u�;�4�Wǿ�&����Q��_�U���;�_�u�u�w�}�W���Y���F��h��3����:�
�
�2��N���DӇ��P	��C1��@��_�u�u�u�w�}�W���Y����Z ��N��U���u�u�0�1�>�f�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�d�h�6������Ƣ�GN��h��*���
�d�|�|�#�8�}���Y���F�N�����7�:��'�"��N������� T��S�����:�9�'��#�i�(߁�����9��d��U���u�u�u�u�w�<��������|��W��E���2�g�b�u�j�<��������|��W������3�
�e�n�-�_������\F��UךU���u�u�u�u�w�}��������A)��hZ��Dۊ�0�
�f�b�k�}��������A)��hZ�����
�
� �d�`��D��Y����G	�G�U���u�u�u�u�w�}��������A��C1�*���'�2�g�m�w�`��������A��C1�*���%��3�
�g�d����Kӂ��]��\����u�u�u�u�w�}�W���&����r��B��L��
�0�
�f�`�a�W���&����r��B��L���8�
�
� �f�j�(��H�ƨ�D��_�N���u�u�u�u�w�}�WϿ�����_'��x��Aӊ�a�'�2�g�n�}�JϿ�����_'��x��Aӊ�0�%��3��m�N���Q����\��XN�\�ߊu�u�u�u�w�}�W�������\
��E!��*���d�
�0�
�d�j�K�������\
��E!��*���!�8�
�
�"�l�@ց�J����W	��C��@��u�u�u�u�w�}�W�������\	��E����
�
�0�
�d�j�K�������\
��E!��*���!�8�
�
�"�l�@ց�J����\��XN�N���u�u�u�u�w�}�WϿ�����_'��x��Aӊ�
�0�
�f�e�a�W���&����r��B��L���8�
�
� �f�j�(��Kӂ��]��G�U���u�u�u�u�w�}��������A��C1�*ي�0�
�f�b�k�}��������A)��hZ�����
�
� �d�`��D������\F��d��U���u�u�u�u�w�<��������|��W��*���
�f�g�i�w�/�(�������F��1�����
� �d�b��n�CϺ�����O��N��U���u�u�u�u�6�/����8����G9��h[�����f�b�i�u�%���������lR��C��*��� �d�b�
�d�h��������l�N��U���u�u�u�4�%�?��������_��h��*��g�i�u�'��2����6����
9��Z��*���d�b�
�f�a�9� ���Y����F�N��U���u�u�4�'�5�2�6�������lQ��R	��F��i�u�'�
�8�1��������G��h8�� ��b�
�f�b�3�*����P���F�N��U���u�4�'�7�8�����&�ߓ�l��h\�G��u�'�
�:�;�/�8���Mʹ��^��h��D��
�f�m�1� �)�W���s���F�N��U���4�'�7�:��/����@�ߓ�V��X�I���'�
�:�9�%����&����l0��B1�Bӊ�f�l�1�"�#�}�^�ԜY���F�N��Uʴ�'�7�:��%�(�(���I����lT��N�U���
�:�9�'��)�Bށ�&����^��G_�U���u�u�u�u�w�}��������A��C1�*���'�2�g�l�w�`����<����|��W�� ��b�
�f�d�w�2����H����F�N��U���u�u�4�'�5�2�6�������lW��E��G��u�h� �
���#���&�ߓ�F9�� _��F��u�:�;�:�f�t�}���Y���F�N�����7�:��'�"��F��&����U��R�� ������ ��d����I�ד� N��
�����d�|�_�u�w�}�W���Y���R��U��4��� �
�d�d��8�(��N���F1��r"��!���
�l�3�
�g�l����Jӂ��]��]����u�u�u�u�w�}�W���&����r��B��D��
�0�
�f�e�a�W���*����g)��h[�����e�d�%�}�c�9� ���Y���9F�N��U���u�u�u�'��2����6����9��h��*��b�i�u����4�������U��Y�����`�1�"�!�w�h�L���Y���F�N��U���
�:�9�'��)�Bށ�&����T��R�� ������ ��d����I�ד� N��S�����|�_�u�u�w�}�W���Y�ƭ�A9��X�����
�d�g�'�0�o�B���Dӓ��`#��t:�����
� �d�b��n�EϺ�����O��N��U���u�u�u�u�6�/����8����G9��h]�����g�b�i�u� ��;���6����
9��h_�D���}�u�:�;�8�n�L���Y���F�N��U���
�:�9�'��)�Bށ�&����T��R�� ������ ��d����I�ד� N��S�����|�_�u�u�w�}�W���Y�ƭ�A9��X�����
�d�`�'�0�o�A���Dӓ��`#��t:�����
� �d�b��n�BϺ�����O��N��U���u�u�u�u�6�/����8����G9��hX�����g�g�i�u� ��;���6����
9��h_�D���}�u�:�;�8�k�L���Y���F�N��U���
�:�9�'��)�Bށ�&����T��R�� ������ ��d����I�ד� N��S�����|�_�u�u�w�}�W���Y�ƭ�A9��X�����
�d�m�'�0�o�O���Dӓ��`#��t:�����
� �d�b��n�OϺ�����O��N��U���u�u�u�u�6�/����8����G9��hW�����g�b�i�u� ��;���6����
9��h_�D���}�u�:�;�8�d�L���Y���F�N��U���
�:�9�'��)�B܁�&����W��R�����7�:��'�"��D�������9��d��U���u�u�u�u�w�<��������|��]��E���2�g�d�u�j�-�F�������]��R
�����2�d�u�:�9�2�F���s���F�N��U���4�'�7�:��/����J����A��\�U��%�d��8�#���������@��_�����:�d�|�_�w�}�W���Y���F��E1�����'� �
�f�f�����K���F��1������4�9�1�>�����Kӂ��]��\����u�u�u�u�w�}�W���&����r��B��F��
�0�
�g�`�a�W���&����G��V�����
�<�}�f�3�*����J��ƹF�N��U���u�u�'�
�8�1��������R��R	��G��i�u�
�
�>�4��������Z��^	��Aʱ�"�!�u�a�l�}�W���Y���F���*���9�'��!�b��B�������F���*���<�<�;�7�2���������W	��C��@��u�u�u�u�w�}�W�������\	��E�����
�
�0�
�f�j�K���&¹��^��r �����<�
�<�}�w�2����H��ƹF�N��U���u�u�'�
�8�1��������9��P1�B���h�%�d��:�)�2�������]9��PF����!�u�|�_�w�}�W���Y���F��E1�����'� �
�f�d�/���N�����h"�����;�7�0�
�9�.�������\F��d��U���u�u�u�u�w�<��������|��]��*���
�d�g�i�w��(�������R��S1��*���}�u�:�;�8�i�L���Y���F�N��U���
�:�9�'��)�B܁�&����W��R������8�!��6�1����&����F��@ ��U���_�u�u�u�w�}�W���Y����Q	��v�� ���f�c�'�2�e�d�W��	�ד�Z��^+�����
�;�&�2�a�9� ���Y����F�N��U���u�u�4�'�5�2�6�������lQ��R	��D��i�u�
�
�>�4��������Z��^	��U���;�:�b�n�w�}�W���Y���F��E�����'��!�`������K���F��1������4�9�1�>�����Y����G	�UךU���u�u�u�u�w�}��������A)��h[��L���2�g�e�u�j�-�F�������]��R
�����2�l�1�"�#�}�^�ԜY���F�N��Uʷ�:�
������������F���G���0�'�<�<��8��������lU��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��G1�����9�d�e�h�2�4����N����U��h�U���u�!�%�3��n�@���Y�ƭ�l��D��ފ�|�|�!�0�]�}�W���Y���F�V�����:�
�:�%�e��B��&����V�
N�����
�:�
�:�'�o�(߁�����9��d��U���u�u�u�u�w�<����&����	��h\��Dߊ�e�3�
�f�w�`��������A9��X��L���3�
�f�d�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2����¹��F��^�����3�
�f�`�'�t����Q����U��Z�����u�%�6�;�#�1�C���P�Ƹ�VǻN��U���u�u�u�u�%���������C9��h_��Dۊ� �g�a�i�w�/�(���?����\	��Y��*���d�b�
�g�]�}�W���Y���F�V�����:�
�:�%�e��B��&���� ^�
N�����
�:�
�:�'�o�(߁�����9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���
�u�u�-�#�2�؁�����9��N�����8�
� �d�c��F������]��[��6���u�=�;�u�w�}�W���Y�����h��3����:�
�b�f��E���&����[��E�����'��:�
�`�m����J�ӓ�]ǻN��U���u�u�u�u�%���������C9��h_��D؊� �f�g�i�w�/�(���?����\	��W��*���d�m�
�g�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʴ�1�}�%�6�9�)����I����K��X ��*���d�f�
�g�w�3�WǪ�	����U��h�Hʴ�
�:�&�
�!��^�������F�N��U���u�u�4�'�;���������9��h_�����m�u�h�4�%�1�(���&����lT��1��*��`�%�n�u�w�}�W���Y�����h��3����:�
�l�f��D���&����[��E�����'��:�
�n�m����J�ד�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Yۇ��P	��C1��D��h�0�<�6�9�j����J�ӓ�O��Y
�����3�
�f�b�'�}�W�������l
��h+��\ʡ�0�_�u�u�w�}�W���Y�ƭ�A9��h(��*���%�g�
�`�f����O���R��[�����:�%�g�
��(�F��&����F�N��U���u�u�4�'�;���������
9��h_�����`�u�h�4�%�1�(���&����lT��1��*��d�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��+�(���Y����P	�� 1��*��`�%�|�4�3�3��������lW�� 1��U���%�6�;�!�;�i�2�������\�C�����f�b�%�u�w�-��������l"���U���}�!�%�3��n�@���Y�ƭ�l��D��ފ�|�u�;�u�8�u��������Q��N�����:�&�
�#��t�W���Y������h��D��
�d�h�4��2����ǹ��F��SN�����8�
� �d�c��F������]��[��L���4�1�;�!��0�(���H����CW������!�9�a�m�~�<�ϰ��θ�C9��h_�B���u�u�%�6�9�)����N����]��X�����3�
�f�b�'�}�W�������l
��hX��U���u�:�}�!�'�;�(��N����F��h�����#�
�|�u�9�}��������F9��Y��D��4�
�:�&��+�(���Y����]	����*���d�a�
�d�j�<�(���
����9��N��ʻ�!�}�8�
�"�l�C؁�H����C9��Y�����g�|�4�1�9�)�_���&���� R��G_��U���6�;�!�9�c�l�^Ͽ�ӈ��N��G1��*��b�%�u�u�'�>�����ғ�O������u�u�u�u�w�}�WϿ�����u	��{��*���d�
�`�3��d�W������G9��E1�����b�e�3�
�d�h���Y���F�N��U���'�
�!��%�����@����S��B1�A��u�'�
�!��/�;���&�ߓ�l ��]�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�d�g�`��������l ��]�*��u�;�u�!�'�;�(��N����F��h�����#�
�|�|�#�8�}���Y���F�N�����9�
�:�
�8�-�E؁�L�ד�F9��N�U���
�!��'��2�(���I����U��h����u�u�u�u�w�}�W���&����\��X��Gӊ�`�f�3�
�g�}�JϿ�����u	��{��*���e�3�
�f�f�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�u�;�u�6�����&����F�R�����b�3�
�f�b�-�^Ͽ��θ�C9��h_�B���u�u�%�6�9�)����K���G��=N��U���u�u�u�u�w�/�(���?����\	��Y��@���3�
�f�u�j�<����&����	��h\��E���
�f�`�%�l�}�W���Y���F���*����'��:��d�Fځ�&����T�
N�����
�:�
�:�'�o�(߁�����9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���
�u�u�-�#�2�؁�����9��N�����8�
� �d�c��F������]��[��D���u�=�;�u�w�}�W���Y�����h��3����:�
�b�f��(���K���F��E1��*���
�:�%�g�����Nƹ��l�N��U���u�u�u�4�%�1�(���&����lT��[��*���g�m�i�u�%���������C9��h^�� ��m�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h_�����}�%�6�;�#�1�F��DӃ��G��SY�� ��f�
�g�u�9�}��������Q��N�����:�&�
�#��t�^Ϫ����F�N��U���u�4�'�9��2�(���	����S��h��G��i�u�'�
�#���������lV��B1�Bߊ�g�_�u�u�w�}�W���Y�ƭ�A9��h(��*���%�g�
�`�1��N���DӇ��l
��q��9���
�l�e�3��n�F���B���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������A	��D�X�ߊu�u�'�6�$�}������ƹF��R	�����u�u�u�3��-���������������h�r�r�u�?�3�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�d�u�9�}��������_��N�����6�;�b�3��n�B���PӇ��N��G1��*��b�%�u�u�'�>�����ғ�O�C�����u�u�u�u�w�}�W���&����\��X��G݊�`�`�3�
�b�}�JϿ�����u	��{��*���e�3�
�f�b�-�L���Y���F�N��U���
�!��'��2�(���Hƹ��U��Z��Hʴ�'�9�
�:��2���&ù��lW��1��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F������%�:�0�&�w�p�W���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�#�
�u�w�%����Ĺ��lW��1��\ʴ�1�}�8�
�"�l�C؁�H����C9��Y�����c�|�u�=�9�}�W���Y���F���*����'��:��j�Fځ�&����R�
N�����
�:�
�:�'�o�(߁�����9��d��U���u�u�u�u�w�<����&����	��h\��Dߊ�
� �f�m�k�}��������l*��G1�*ڊ� �d�m�
�e�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3����H�����C��݊� �d�f�
�e�}��������F9��Y��D��4�
�:�&��+�(���PӒ��]l�N��U���u�u�u�4�%�1�(���&����lT��[��*���g�m�i�u�%���������C9��h^�� ��b�
�g�_�w�}�W���Y���F��E1��*���
�:�%�g��h�@���&����[��E�����'��:�
�n�m����J�ד�]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Yۇ��P	��C1��D��h�0�<�6�9�j����J�ӓ�O��Y
�����3�
�f�b�'�}�W�������l
��hV��\ʡ�0�_�u�u�w�}�W���Y�ƭ�A9��h(��*���%�g�
�`�o�;�(��Y����A��C1�����:�
�b�e�1��D���	��ƹF�N��U���u�u�'�
�#���������lW��1��*��u�h�4�'�;���������
9��Q��F���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U´�
�:�&�
�!��W�������]��Q��F���%�|�4�1��0�(���H����CW������!�9�a�l�~�}����Y���F�N��U���'�
�!��%�����N����
9��h\�U��4�'�9�
�8�����KĹ��U��Y����u�u�u�u�w�}�W�������G9��E1�����l�d�
�
�"�n�G��Y����_��X�����g�
�
� �f�e�(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�4�3�u��������EW��S�����:�1�
� �f�n�(��Y������h��D��
�d�h�4��2����ǹ��O��_��U���u�u�u�u�w�}��������A9��X��B��
� �g�e�k�}��������l*��G1�*ڊ� �d�b�
�e�W�W���Y���F�N�����
�:�
�:�'�o�(���M���� W��S�����!��'��8��N�������W��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��RN�����!�!�u�4������Y����[��C��U���=�;�{�x�]�}�W���7����^9��D��*���6�o�%�:�2�.�_���:����^J��G1��Yʴ�
�<�
�1��l�[ϻ�����WQ��B1�Fߊ�g�_�u�u�2�4�}���Y���P����6���&�u�&�u�w�}�W���Yӑ��]F��h=�����3�8�e�h�w�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����4�
�<�
�3��F���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=�����3�8�d�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����3�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]´�
�:�&�
�!��W�������]��Q��F���%�|�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��h^�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�)����D���F�N��U���u�u�4�
��;���YѾ��l�N��Uʰ�1�6�&�n�w�}����	����@��=N��U���4�
�:�0�6�.��������@H�d��Uʴ�
�:�0�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��B�����:�1�
� �f�n�(��s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ����F��*���&�
�#�
�w�}��������U��]�����|�u�=�;�]�}�W���Y���R��X ��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������_��D��ʥ�:�0�&�u�z�}�WϿ�&����l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��^���Yӄ��ZǻN��U���3�}�;�!��-��������Z��S�����4�!�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�<�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�%�<�Ͽ�
����C��R��U���u�u�4�
�2�9�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����y�0�<�6�9�j����J�ӓ�OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���K����lW�V �����}�%�6�;�#�1�F��DӃ��G��SY�� ��f�
�g�|�~�)����Y���F�N�����4�,�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��A��NN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����1�
�e�u�$�4�Ϯ�����F�=N��U���&�2�7�1�f�m��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e��.����8����R��[
��U���7�2�;�u�w�}�W���Y�����D�����d�e�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��Y������b�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��D�����
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����I���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�e� �$�<����&˹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����d�m�4�&�0�}����
���l�N��*���
�1�
�d��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�;�4�1����@����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����f��V��4���
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����K�ƭ�@�������{�x�_�u�w�-��������Q��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�]��[��<��
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e� �&�6�8�6���I����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����f�u�&�<�9�-����
���9F������7�1�d�c�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�e� �&�6�8�6���H����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����f��V��4���d�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����H����R��P �����&�{�x�_�w�}��������lW��1�����
�'�6�o�'�2��������T9��R��!���g�3�8�d�w�%����Ĺ��lW��1��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�b�u�j�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�#��}�W�������9��h_�@���|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�d�W�������A	��D�X�ߊu�u�%�&�0�?���@ù��@��h����%�:�0�&�#�-����J�ѓ�OǻN�����_�u�u�u�w�}�W���Y����Z��S
��F��i�u�;�!��0�(���H����CW������!�9�a��~�<�ϰ��θ�C9��h_�B���u�u�%�6�9�)����=����]��X�����3�
�f�b�'�}�W�������l
��h-��U���u�:�}�!�'�;�(��N����F��h�����#�
�|�u�9�}��������F9��Y��D��4�
�:�&��+�(���Y����]	����*���d�a�
�d�j�<�(���
����9��N��ʻ�!�}�8�
�"�l�C؁�H����C9��Y�����m�|�4�1�9�)�_���&���� R��G_��U���6�;�!�9�c�j�^Ͽ�ӈ��N��G1��*��b�%�u�u�'�>�����ғ�O��Y
�����!�%�3�
�d�j����Y����\��h��*���u�;�u�:��)����&����l��
N��*���&�
�#�
�~�}��������^��B1�A݊�d�h�4�
�8�.�(���&���R��Y��]���
� �d�a��l�JϿ�&����G9��1�\ʴ�1�;�!�}�:����MĹ��[��G1�����9�a�d�|�6�9����Q����U��Z�����u�%�6�;�#�1�C��P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��[�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�� ���4�0��
�e�<�(���P�����^ ךU���u�u�u�u�w�}��������lW��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������r/��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�i�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(�������r/��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�c�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���6�9�1��f���������F�R �����0�&�_�_�w�}�ZϿ�&����Q��X����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���6�9�1��f��������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�G���
����W'��Z�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��j�W�������A	��D�X�ߊu�u�%�&�0�?���K����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�G���
����W'��[�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�`�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��E���&�4�0���h�������9F���U���6�&�n�_�w�}�Z���	����l��h_����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�d�u�j�u����&����F��@ ��U���h�4�
�:�$��ށ�P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Mۊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��h_�����<�;�7�0��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����^��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�l�;�������Q
��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�n�}����Ӗ��P��N����u�%�&�2�5�9�F�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�h�?���5����lV��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�l�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����8�!�e�4��1�^��Y����]��E����_�u�u�x�w�-��������
_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9����9���!�d�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����H���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�>�5����&¹��l��G�U���0�1�%�:�2�.�}�ԜY�����D�����g�m�4�&�0�}����
���l�N��*���
�1�
�e��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�<�?�4����&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��G��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ӓ�Z��^��*؊�%�#�1�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�L����[*��^��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��l�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������2��8�#�n�������9F���U���6�&�n�_�w�}�Z���	����l��h\�U���<�;�%�:�2�.�W��Y����C9��P1����c�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��@���2��8�!�c�<�(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������G9��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�b�<����Y����V��C�U���4�
�<�
�3��Dځ�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u����������9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�g�`�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h&�����<�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Z�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lS��^	�����
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����M���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�`��0�����O����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����`�u�&�<�9�-����
���9F������7�1�g�f�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�`��2��0��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��@���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&ƹ��T��Z��B���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&������C1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�e�o�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ߊ�<�=�<�<����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��Y����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���=�<�<�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����Q��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�h�?���5����l_��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�m�w�.����	����@�CךU���%�&�2�7�3�o�G���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�b���������9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�g�e�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h&�����<�
�e�4��1�^��Y����]��E����_�u�u�x�w�-��������_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��V�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9����9���!�d�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�`��:�;�������R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�g�m�4�$�:�W�������K��N�����<�
�1�
�n���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�>�5����&�ԓ�C9��SGךU���0�<�_�u�w�}�W���Y���R��^	�����l�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��P�����d�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lU��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l.��_"�����f�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���N�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�<�?�4����J����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����d�u�&�<�9�-����
���9F������7�1�f�c�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�`��2��0���&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��F��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ӓ�Z��^��*���4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���LӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ƹ��T��Z��Dߊ�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��E���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`��2��:�)�Fځ�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��F��4�&�2�u�%�>���T���F��h��*���
�f�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���
�:��8�#�m������ƹF��R	�����u�u�u�u�w�}�W���
����W��Z��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�����Z��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�c�}����Ӗ��P��N����u�%�&�2�5�9�D�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�j�;�������9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�f�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h"��9���!�d�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��@"�����
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�b��"�>�4�(݁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��F��4�&�2�u�%�>���T���F��h��*���
�c�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���
�:��8�#�n������ƹF��R	�����u�u�u�u�w�}�W���
����W��_��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(؁�����Z��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�`�<����Y����V��C�U���4�
�<�
�3��@���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�g���������9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�u�h��<�(���
����T��N����� �&�4�0���(������R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W�� ^�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lQ��X�����a�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���I�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�:��0��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�l�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b��"�<�>��(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Y�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����5����^��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�d�e�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(���5����lP��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F�� 1�����<�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Y�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lQ��X�����b�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���N�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�:��0��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�c�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b��"�<�>��(������F�U�����u�u�u�u�w�}�WϿ�&����Q��^�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����5����^��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�c�h�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(���5����l_��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�d�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F�� 1�����<�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Z�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lQ��X�����d�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����K���N��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b�� �4����I����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����f�u�&�<�9�-����
���9F������7�1�a�f�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�b��"�>�4�(�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��F���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��D*��^��D���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����Z��h_�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�o�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*݊�:��8�!�f���������F�R �����0�&�_�_�w�}�ZϿ�&����Q��[����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*����8�!�d��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����S��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�;�������U��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�6�.��������@H�d��Uʴ�
�<�
�1��k��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e��.����8����R��[
��U���7�2�;�u�w�}�W���Y�����D�����a�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��D�����
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lR��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l*��{����
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��Y���]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�b��"�>�4�(�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�a�l�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b��"�<�>��B���&����9F����ߊu�u�u�u�w�}�W���	����l��hZ�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����Z��h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�i�GϿ�
����C��R��U���u�u�4�
�>�����Aù��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ց�����V��Z�����;�4�
�9�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���I�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�;�4�1��������[/��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�a�f�<����Y����V��C�U���4�
�<�
�3��Nށ�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u��l�"�������Z��{�����
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�i�F��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���d� �&�4�2���������R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�`�e�4�$�:�W�������K��N�����<�
�1�
�g���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�g��8��������l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1�����e�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��9��R�����
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����LӇ��Z��G�����u�x�u�u�6���������l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ϯ�I����P��S/��G���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�h�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N����� �&�4�0���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Aʴ�&�2�u�'�4�.�Y��s���R��^	�����d�
�&�<�9�-����Y����V��V�����y�%�e� �$�<����&ù��l��h�����u�
�
�;�4�1����H����E
��^ �����%�e� �&�6�8�6���&����_��Y1�����
�
�;�6�;�9�>�������W9��h��Yʥ�e� �&�4�2��(ہ�	����l��D��U���
�;�6�9�3��B���&����Z��^	���� �&�4�0���(�������]9��PB��*ڊ�;�6�9�1��j��������l��N��E���&�4�0�����������@����*���6�9�1��n�<�(���&����Z�G1�� ���4�0��
�g�<�(���&����Z�G1�� ���4�0��
�f�<�(���&����Z�G1�� ���4�0��
�e�<�(���&����Z�G1�� ���4�0��
�d�<�(���&����Z�G1�� ���4�0��
�c�<�(���&����Z�G1�� ���4�0��
�b�<�(���&����Z�G1��9���!��4�9�3�<�(���&����Z�G1��=����8�!�e�6���������F��1�����8�!�d�4��1�(���
���C9����9���!�g�4�
�;������Ƽ�9��P�����f�4�
�9��3����Y����{��{�����4�
�9�
�9�.����&ƹ��T��Z��@���
�9�
�;�$�:�W���&������C1�����9�
�;�&�0�}�(ځ�����^�� 1��*���
�;�&�2�w��(�������G9��V�����;�&�2�u����������
9��h��*���&�2�u�
��4��������l��A�����<�y�%�`��:�;�������R��[
�����2�u�
�
�>�5����&�ԓ�C9��S1��*���y�%�`��0�����H����l��h�����u�
�
�<�?�4����M����E
��^ �����%�`��2��0���&����_��Y1�����
�
�:��:�)�G���&����Z��^	�����"�<�<����������@����*����8�!�g�6���������F�� 1�����<�
�
�%�!�9��������lQ��X�����a�4�
�9��3����Y����	��^��*ߊ�%�#�1�<��4�[Ϯ�N������C1�����9�
�;�&�0�}�(؁�����Z��h�����<�
�<�y�'�j�;�������9��h��*���&�2�u�
��2�;����ߓ�C9��S1��*���y�%�b�� �4����I����E
��^ �����%�b��"�>�4�(�������W9��h��Yʥ�b��"�<�>��E���&����Z��^	�����"�<�<��n��������l��N��B���"�<�<�
�c�<�(���&����Z�G1��9���<�<�
�`�6���������F��1�����0��8�!�>�5����&����Z��^	���
�;�6�9�3�4��������C9��S1��*���y�%�d�
�;�<�;�������E
��^ �����u�u�7�2�9�}�W���Y���F������7�1�c�a�k�}�_���K����R��Z�����9�
�;�&�0�`��������_	��T1�U���}�
�d� �$�<��������D/��V�����;�&�2�h�6�����&����P9����]���
�;�6�9�3�4��������R��[
�����2�h�4�
�8�.�(�������	����*���<�<�;�7�2���������@��
N��*���&�
�:�<��t����	�ӓ�Z��^��*ڊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`��:�;����ד�C9��S1��*���u�u�%�6�9�)�������\�G1��=����8�!�g�6���������[��G1�����9�2�6�e�w�/�_���&������C1�����9�
�;�&�0�`��������_	��T1�U���}�
�
�<�?�4����&����_��Y1����4�
�:�&��2����PӉ����h&�����<�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�B�������Z��h�����<�
�<�u�w�-��������Z��N��U¥�`��2��:�)�@���&����Z��^	��U���6�;�!�9�0�>�G����μ�9��P�����m�4�
�9��3����DӇ��P	��C1�����e�u�'�}����������
9��h��*���&�2�h�4��2��������O��EN��*ߊ�<�=�<�<��m��������l��S�����;�!�9�2�4�m�W���Q����{��{����
�%�#�1�>�����Y����\��h�����|�:�u�%�b���������9��h��*���&�2�h�4��2��������O��EN��*ߊ�<�=�<�<��n��������l��S�����;�!�9�2�4�m�W���Q����{��{����
�%�#�1�>�����Y����\��h�����|�:�u�%�b���������9��h��*���&�2�h�4��2��������O��EN��*݊�:��8�!�g�<�(���&����Z������!�9�2�6�g�}����&Ĺ��D*��^��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�b�� �4����&����_��Y1����4�
�:�&��2����PӉ����h"��9���!�f�4�
�;���������C9��Y�����6�e�u�'���(���5����lR��G1�����
�<�u�u�'�>��������lV�X������"�<�<����������@��
N��*���&�
�:�<��t����	�ѓ�\��Z��C���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�8�����N����E
��^ �����u�%�6�;�#�1����I�ƣ�N�� 1�����<�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�@�������G9��V�����;�&�2�h�6�����&����P9����]���
�:��8�#�l�(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l*��{����
�%�#�1�>�����Y����\��h�����|�:�u�%�`�� �������l��A�����<�u�u�%�4�3��������F��F��B���"�<�<�
�d�<�(���&����Z������!�9�2�6�g�}����&Ĺ��D*��^��A���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�8�����Hƹ��l��h�����h�4�
�:�$�����&����AF��h^�����9�1��e�6���������[��G1�����9�2�6�e�w�/�_���&����R
��v'��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�e� �$�<����&����l��h�����h�4�
�:�$�����&����AF��h^�����9�1��f�6���������[��G1�����9�2�6�e�w�/�_���&����R
��v'��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�e� �$�<����&ƹ��l��h�����h�4�
�:�$�����&����AF��h^�����9�1��c�6���������[��G1�����9�2�6�e�w�/�_���&����R
��v'��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�e� �$�<����&˹��l��h�����h�4�
�:�$�����&����AF��h^�����9�1��l�6���������[��G1�����9�2�6�e�w�/�_���&����R
��v'��E���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�9�>����0����R��[
�����2�h�4�
�8�.�(�������	����*���6�9�1��f���������@��
N��*���&�
�:�<��t����	�֓�]��[��<��
�%�#�1�>�����Y����\��h�����|�:�u�%�g���������R��G1�����
�<�u�u�'�>��������lV�X����� �&�4�0���B���&����Z��^	��U���6�;�!�9�0�>�G����έ�l��E��U���6�;�!�9�0�>�G���s���V��G�����_�_�u�u�z�<�(���&����W��V�����'�6�&�{�z�W�W���	����l��hX�*���<�;�%�:�w�}����
�έ�l��h�����
�!�
�&��q��������W9��GךU���0�<�_�u�w�}�W���Y���R��^	�����d�u�h�}�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����2�7�1�c�c�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����R��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�]��[��<���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�A���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�e� �&�4�2��(܁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��B���&�<�;�%�8�8����T�����D�����b�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ڊ�;�6�9�1��i������ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�G���
����W'��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�k�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����W��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�}����Ӗ��P��N����u�%�&�2�5�9�O݁�
����l��TN����0�&�4�
�#�/�[Ͽ�&����P��h=�����3�8�e�u����������lS��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�g�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h;�����1��`�4��1�^��Y����]��E����_�u�u�x�w�-��������F��D��U���6�&�{�x�]�}�W���
����W��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��D�����
�
�%�#�3�W�W�������F�N��U���u�u�4�
�>�����H�����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�;�4�1����O����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����`�u�&�<�9�-����
���9F������7�1�l�a�6�.���������T��]���&�2�6�0��	��������F��^�����3�
�f�`�'�t�W�������9F�N��U���u�u�u�%�$�:����@���F�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1�9�)�_�������l
��h^��U���!�:�1�
�"�l�Dځ�K���9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lW��=N��U���<�_�u�u�w�}����	����l��h_�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�o����H����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���
����@��d:��؊�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�'��2����6����
9��Q��G���%�u�h�4�%�?��������_��R��#���
�e�l�%��}�W�������V�=N��U���
�:�9�'��)�Cց�����l ��^�*��i�u�u�u�w�}��������_��h^�����}�:�9�-�����&����P��G\��\��r�r�u�9�2�W�W���Y�Ƽ�
9��D�����8�!�<�=�9�4�(���B�����h������!�`�
��(�F��&���F��h=��0��� �
�l�3��m�F���Q���F��@ ��U���_�u�u�'��2����6���� 9��Q��Fߊ�d�i�u�
��4��������W9��h��]���u�u�:�;�8�m�L���YӇ��l
��q��9���
�b�e�3��n�B���Y���Q	��h �����'�
�a�3��n�D���Y����Q	��h��3����:�
�c�'�4����@ù��O��N�����9�
�:�
�8�-�Eց�&���� ^��G\��H���:�9�;�1��8���&���� P��G\�����:�9�9�
�8�����KŹ��Z9��hV�*��|�_�u�u�z�}��������A9��X��G���<�3�
�d��n�W�������A	��D�X�ߊu�u�:�9�;���������9��^1��*��
�f�
�&�>�3����Y�Ƽ�\��DF�����:��'� ��d�G�������J��E�����'��!�a������J���R��U��4��� �
�l�g�%�:�E��UӇ��l��[/��:���a�
�
�0��n�@�������\
��E!��*���a�'�2�g�c�q��������A��C1�*ߊ�0�
�f�b�w�/�(�������F��1�����g�`�y�4�%�?��������_��h��*��b�u�'�
�8�1��������9��P1�C���4�'�7�:��/����@�ߓ�V��X�U���
�:�9�'��)�Cց�I����lT��B�����:�9�'��#�i�(������� Q����*���9�'��!�c��E�������J��E�����'��!�a��n����K������h������!�a�
�c�/���@����A��X�����!�a�
�`�%�:�E��UӒ��l ��]�*��u�%�&�2�5�9�F��UӇ��@��U
��D��|�u�u�7�0�3�W���Y����UF��G1�����1�d�b�|�#�8�}���Y���F�^��]���
� �d�a��l�JϿ�&����G9��1�\ʡ�0�u�u�u�w�}�W���Y����\	��[�����:�%�g�
�?����O����Z�V������'� �
�n�m����K����9F�N��U���u�9�<�u�6���������
V�C��U���u�u�u�u�w�}�Wϼ�����l ��h"����
�=�
� �o�k���E�ƭ�A9��X�����
�l�d�
�2��D��s���F�N�����3�}�!�%�1��D���	���R��X ��*���
�|�u�=�9�W�W���Y���F�N�����!��'��8��E�������W��G]�I���'�
�:�9�%����&�ғ�V��W����u�u�u�u�w�1����Q����U��Z�����u�%�6�;�#�1�C���PӒ��]FǻN��U���u�u�u�u�8�1��������\��1�����
�d�
�f�w�`��������A��C1�*���'�2�g�m�l�}�W���Y�����^��]���
� �d�a��l�JϿ�&����G9��1��\ʡ�0�u�u�u�w�}�W���Y����\	��[�����:�%�g�
�?����O����Z�V������'� �
�n�l�(���&����l�N��U���u�0�&�3��)����&����l��
N��*���&�
�#�
�~�}����s���F�N��U���7�:�
�!��/�;���&�ԓ�[��B1�C���g�i�u�'��2����6����
9��h��*��b�_�u�u�w�}�W�������N��G1��*��b�%�u�u�'�>�����ғ�O��_�����u�u�u�u�w�}�W�������u	��{��*���%�<�3�
�f��D���DӇ��l��[/��:���a�
�e�'�0�o�@��Y���F�N�����u�}�8�
�"�l�C؁�H����C9��Y�����l�|�!�0�w�}�W���Y���F������
�:�
�:�'�o�(���&����P��\��Hʴ�'�7�:��%�(�(���@����lT�� UךU���u�u�u�u�;�4�W�������lW�� 1��U���%�6�;�!�;�i�O�������9F�N��U���u�u�u�:�;�1�(���&����lT��G�����d�
�f�u�j�<��������|��W��*���
�f�g�_�w�}�W���Y�Ʃ�@��F�����
�f�b�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����l
��q��9���
�g�%�<�1��Fف�J�����h������!�a�
��8�(��N���F�N��Uʰ�&�3�}�!�'�;�(��N����F��h�����#�
�|�u�?�3�}���Y���F�N�����
�!��'��2�(���	����F9��1��G��u�'�
�:�;�/�8���Mʹ��A��]�N���u�u�u�u�w�8����Qے��l ��]�*��h�4�
�:�$��ہ�P�Ƹ�V�N��U���u�u�u�u�5�2�(���?����\	��\����� �m�c�%�e�a�W���&����r��B��L���'�2�g�a�l�}�W���Y�����^��]���
� �d�a��l�JϿ�&����G9��1�\ʡ�0�u�u�u�w�}�W���Y����\	��[�����:�%�g�
�?����O����Z�V������'� �
�n�i����K����9F�N��U���u�9�<�u��0�(���H����CW������!�9�a�f�~�)����Y���F�N��U���:�9�9�
�8�����K����Z9��hV�*��u�h�4�'�5�2�6�������lU��R	��F��_�u�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}��������A9��X��G���<�3�
�d��n�W������\	��E����
�
�0�
�d�o�}���Y���F�R�����!�%�3�
�d�j����Y����\��h��*���u�=�;�_�w�}�W���Y���F��X�����'��:�
�e�-����&����CU��S�����:�9�'��#�i�(ށ�����Q��N��U���u�u�0�&�w�}�W���Y���F������
�:�
�:�'�o�(���&����P��\��H���w�_�u�u�w�}�W����ƥ�l�N��Uʰ�&�u�u�u�w�}�W�������_��X�����g�
�=�
�"�e�A���K���>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�:�9�;���������9��^1��*���
�f�u�&�>�3�������KǻN�����9�
�:�
�8�-�Eہ�����l^��h�*���<�;�%�:�w�}����
�έ�A9��X�����
�d�e�'�0�o�C������\	��E�����
�
�0�
�e�j�W���&����r��B��D���'�2�g�`�{�<��������|��_��*���
�g�b�u�%���������lS��1����c�y�4�'�5�2�6�������lS��R	��G��u�'�
�:�;�/�8���L¹��A��\�Yʴ�'�7�:��%�(�(���N����lT�� B�����:�9�'��#�h�(ׁ�����T�V������'� �
�f�d����K������h������!�`�
�g�/���@����A��X�����!�`�
�d�%�:�E��UӇ��l��[/��:���`�
�g�'�0�o�G������\	��E�����
�f�'�2�e�m�[Ͽ�����_'��x��@ۊ�a�'�2�g�f�q��������A��C1�*���'�2�g�d�{�)����&����l�������7�1�d�l�{�<�(���&����U��d��Uʷ�2�;�u�u�w�}��������T9��S1�B���!�0�_�u�w�}�W���Y�����h��D��
�d�h�4��2����ǹ��F��R ��U���u�u�u�u�w�}����&����\��X��Gފ�=�
� �m�d�-�E��Y����Q	��v�� ���d�e�'�2�e�i�L���Y���F������4�
�<�
�3��D��Y����l�N��U���u�u�u�7�8���������C9��h��*���m�f�%�g�k�}��������A)��h[��Dߊ�0�
�f�b�]�}�W���Y���V
��QN�����3�
�f�b�'�}�W�������l
��h+��U���;�_�u�u�w�}�W���Y�Ʈ�\
��C1�����:�
�a�%�>�;�(��&����[��E�����'��!�`��i����K����9F�N��U���u�9�<�u��0�(���H����CW������!�9�a��~�)����Y���F�N��U���:�9�9�
�8�����Kǹ��Z9��hV�*��u�h�4�'�5�2�6�������lW��E��G��n�u�u�u�w�}�Wϻ�
�����h��D��
�d�h�4��2����ǹ��F��R ��U���u�u�u�u�w�}����&����\��X��Gފ�=�
� �m�d�-�E��Y����Q	��v�� ���d�d�
�0��n�E�ԜY���F�N�����}�!�%�3��n�@���Y�ƭ�l��D��ފ�|�u�=�;�]�}�W���Y���F�U��*����'��:��i�������� 9��N�U���
�:�9�'��)�Bށ�H����lT�� UךU���u�u�u�u�;�4�W�������lW�� 1��U���%�6�;�!�;�i�6�������9F�N��U���u�u�u�:�;�1�(���&����lT��G�����`�
�f�u�j�<��������|��_��E���2�g�l�n�w�}�W���Y����_��F����� �d�a�
�f�`��������_��G�����u�u�u�u�w�}�W���Yӄ��_9��h(��*���%�g�
�=��(�O���	���F��E1�����'� �
�d�n�/���A��ƹF�N��U���9�<�u�}�:����MĹ��[��G1�����9�a�m�|�#�8�W���Y���F�N��U���9�9�
�:��2���&����U��]��F���h�4�'�7�8�����&�ד�l��h\�G�ߊu�u�u�u�w�}����Y�θ�C9��h_�B���u�u�%�6�9�)����N����[��=N��U���u�u�u�u�w�2����&����	��h\�����3�
�`�
�d�}�JϿ�����_'��x��@ۊ�
�0�
�g�`�W�W���Y���F��D��]¡�%�3�
�f�`�-�W���	����@��AZ��\���=�;�_�u�w�}�W���Y���Q	��h��3����:�
�a�'�4����L����F���*���9�'��!�b��(���&����l�N��U���u�0�&�3��)����&����l��
N��*���&�
�#�
�~�}����s���F�N��U���7�:�
�!��/�;���&�ғ�[��B1�F���g�i�u�'��2����6����9��E��G��n�u�u�u�w�}�Wϻ�
�����h��D��
�d�h�4��2����ǹ��F��R ��U���u�u�u�u�w�}����&����\��X��Gފ�=�
� �m�d�-�E��Y����Q	��v�� ���d�a�'�2�e�k�L���Y���F������}�8�
� �f�i�(��DӇ��P	��C1��A��|�!�0�u�w�}�W���Y���F��X�����:�
�:�%�e���������l��R�����7�:��'�"��F�������S��=N��U���u�u�u�9�>�}�_���&���� R��G_��U���6�;�!�9�c�o�^Ϫ���ƹF�N��U���u�u�:�9�;���������9��^1��*���
�f�u�h�6�/����8����G9��h\�����g�g�_�u�w�}�W���Y����UF�C�����f�b�%�u�w�-��������lW����ߊu�u�u�u�w�}�W�������G9��E1�����a�%�<�3��h�(��Y����A��X�����!�`�
�
�2��E��s���F�N�����u�u�u�u�w�}�W���Yӄ��_9��h(��*���%�g�
�=��(�O���	���F��UךU���u�u�u�u�9�}��ԜY���F��D��U���u�u�u�u�5�2�(���?����\	��Z����� �m�f�%�e�a�W͆�B���F���U���u�u�u�0�3�-����
��ƓF�C�����9�
�:�
�8�-�Eف�����l^��h�U���<�;�%�:�2�.�W��Y����\	��[�����:�%�g�
�?����I����l��^	�����u�u�'�6�$�u��������A)��h[��E���2�g�c�y�6�/����8����G9��h_�����d�b�u�'��2����6���� 9��E��G��y�4�'�7�8�����&�Փ�l��h\�B���'�
�:�9�%����&ǹ��T9��\����7�:��'�"��D�������^����*���9�'��!�b��(���&����F��E1�����'� �
�f�`�/���@����A��X�����!�`�
�
�2��E��Y����Q	��v�� ���f�l�'�2�e�m�[Ͽ�����_'��x��@ي�e�'�2�g�f�q��������A��C1�*���'�2�g�d�{�<��������|��]��G���2�g�g�y�6�/����8����G9��h_�����g�g�y�4�%�?��������U��1����f�y�4�'�5�2�6�������lW��E��G��y�!�%�3��n�@���UӇ��@��U
��D��y�4�
�<��9�(��O���F��P��U���u�u�<�u�6���������P�C�����u�u�u�u�w�;�_Ǫ�	����U��h�Hʴ�
�:�&�
�!��^������F�N��U���u�u�7�:��)�1���5����P��_�� ��e�%�g�i�w�/�(�������F��1�����g�c�n�u�w�}�W���YӃ��Z �V�����1�
�f�e�w�5��ԜY���F�N��Uʷ�:�
�!��%�����O����l ��W����i�u�'�
�8�1��������S��R	��G��_�u�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}��������A9��X��C���<�3�
�l��n�W������\	��E�����
�a�'�2�e�n�L���Y���F������}�8�
� �f�i�(��DӇ��P	��C1��A���|�!�0�u�w�}�W���Y���F��X�����:�
�:�%�e���������l��R�����7�:��'�"��D��&����T��d��U���u�u�u�0�$�;�_Ǫ�	����U��h�Hʴ�
�:�&�
�!��^������F�N��U���u�u�7�:��)�1���5����P��_�� ��e�%�g�i�w�/�(�������F��1�*���
�g�g�_�w�}�W���Y�Ʃ�@��F�����
�f�b�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����l
��q��9���
�c�%�<�1��N߁�J�����h������!�`�
�f�/���H��ƹF�N��U���9�<�u�}�:����MĹ��[��G1�����9�a��|�#�8�W���Y���F�N��U���9�9�
�:��2���&����U��^��F���h�4�'�7�8�����&�Փ�9��P1�D��u�u�u�u�w�}��������^��B1�A݊�d�h�4�
�8�.�(���&���G��d��U���u�u�u�u�w�?��������l*��G1�*���
� �m�e�'�o�K�������\
��E!��*���l�'�2�g�g�f�W���Y���F��[��U���8�
� �d�c��F������]��[��M���!�0�u�u�w�}�W���Y�����[1��*���
�:�%�g��5�(���A�֓� T�
N�����:��'� ��n�O�������]ǻN��U���u�u�9�<�w�u��������9��S�����;�!�9�a�`�t����Y���F�N��U���u�:�9�9��2�(���	����C��Q��Lڊ�f�u�h�4�%�?��������U��h��*��b�_�u�u�w�}�W�������N��G1��*��b�%�u�u�'�>�����ғ�O��_�����u�u�u�u�w�}�W�������u	��{��*���%�<�3�
�n��D���DӇ��l��[/��:���`�
�
�0��l�E�ԜY���F�N�����}�!�%�3��n�@���Y�ƭ�l��D��ފ�|�u�=�;�]�}�W���Y���F�U��*����'��:��k��������9��N�U���
�:�9�'��)�B܁�&����W��d��U���u�u�u�0�$�;�_Ǫ�	����U��h�Hʴ�
�:�&�
�!��^������F�N��U���u�u�7�:��)�1���5����P��_�� ��e�%�g�i�w�/�(�������F��1�����g�m�n�u�w�}�W���YӃ��Z ���*���d�a�
�d�j�<�(���
����9��N�����u�u�u�u�w�}�W�������_��X�����g�
�=�
�"�e�G���K���R��U��4��� �
�f�f�%�:�E��B���F�N��U���<�u�}�8��(�F��&�����T�����a�g�|�!�2�}�W���Y���F�N�����9�
�:�
�8�-�Eف�����l^��h�U��4�'�7�:��/����J�ԓ�V��Y����u�u�u�u�w�1����Q����U��Z�����u�%�6�;�#�1�C��PӒ��]FǻN��U���u�u�u�u�8�1��������\��1�����
�l�
�f�w�`��������A��C1�*ۊ�0�
�d�b�]�}�W���Y���V
��d��U���u�u�u�u�w�?��������l*��G1�*���
� �m�e�'�o�K���!��ƹF�N��U���;�u�3�_�w�}�W������F�N��U���7�:�
�!��/�;���&�Г�[��B1�E���g�i�u��l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W�������]	��h����
� �d�c��o�K�������K!��x��Fۊ� �d�`�
�e�2�W�������u	��{��*���%�<�3�
�f��D���s���Q	��h �����'�
�b�3��n�N���Y���Q	��h�����
�c�3�
�d�j����ӄ��_9��h(��*���%�g�
�=��(�O���	���9F��������!�f��(�F��&���F�N�����&�2�0�}� �1�(���&����lW��G�����e�
�f�|�i�.����Q����G9��E1�����m�%�<�3��i�(��P�Ʃ�@�L�U���7�:�
��.�(�(���I����U��[�����h�}�:�9���5�������G9��h^�����%�6�;�!�;�l�F��Y����\	��O)��:���c�
� �d�a��G��Y���C9��h-�����8�!�<�
�>�q�������A�=N��U���9�-���#�k�(���H����CT�
N�����-���!�a����Oƹ�����������!�c��)����&����l��d��Uʷ�:�
��,�"��A���&����l��S��D���=�;�}�<�9�9��������l*��G1�*���
� �b�`�'�o�W���������[�����:�%�g�
�?����@����O��[��W���_�u�u�-�#�2�؁�����9��R��W���"�0�u�<��4�1���5����@9��P1�D��4�
�:�&��+�(��Y����D��d��Uʼ�
�<��'��2�(�������W��N�U���
�:�<�
�2�)�ǫ�
����WN��h��3����:�
�
�2��N���Rӓ��Z��SF��*���&�
�#�
�~�f�}���Y����d9��h(��*���%�d�
�=��(�@���	����@��YN�����&�u�x�u�w�4�(���?����\	��X����� �b�`�%�e�<����&����\��E�����
�
�;�6�;�9�>�������TJ��h^�����9�1��d�>����	�֓�]��[��<���<�
�<�y�'�m�"�������z9��^ �����%�e� �&�6�8�6���&����Z�G1�� ���4�0��
��3����Y����f��V��4���
�;�&�2�w��(�������r/��h�����u�
�
�;�4�1����A����@����*���6�9�1��n�4�(���UӖ��l3��T�����d�
�;�&�0�}�(߁�����V��h_�����<�y�%�e��.����8����l��D��U���
�;�6�9�3��F܁�����F��1�����0��
�a�>����	�֓�]��[��<��
�;�&�2�w�0�(���H����CW�V�����1�
�f�e�w�-�������� Q��=N��U���<�_�u�u�w�}����	����l��h_�C���=�;�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}� ���&����	��h_�����3�
�e�
�d�}�JϮ�I����P��S/��E���
�<�n�u�w�}�W���YӃ��Z �V�����1�
�f�e�w�5��ԜY���F�N��Uʼ�
�!��'��2�(���	����F9��1��G��u�
�
�;�4�1����Hƹ��l��d��U���u�u�u�0�$�;�_Ǫ�	����U��h�Hʴ�
�:�&�
�!��^������F�N��U���u�u�<�
�#���������l��h��B���%�g�i�u����������lW��^ ����u�u�u�u�w�}��������^��B1�A݊�d�h�4�
�8�.�(���&���G��d��U���u�u�u�u�w�4�(���?����\	��X����� �b�`�%�e�a�W���&����R
��v'��F���
�<�n�u�w�}�W���YӃ��Z ���*���d�a�
�d�j�<�(���
����9��N�����u�u�u�u�w�}�W�������l ��h"����
�=�
� �`�h���E�Ƽ�9��D�����
�g�<�
�>�f�W���Y���F��[��U���8�
� �d�c��F������]��[��7���!�0�u�u�w�}�W���Y�����[�����:�%�d�
�?����L����Z�G1�� ���4�0��
�f�4�(���B���F�N��U���<�u�}�8��(�F��&�����T�����a��|�!�2�}�W���Y���F�N��"���
�:�
�:�'�l�(���&����S��\��Hʥ�e� �&�4�2��(�������T]ǻN��U���u�u�9�<�w�u��������9��S�����;�!�9�a�n�t����Y���F�N��U���u��9�
�8�����HŹ��Z9��hY�*��u�h�%�e��.����8����Z��^	�U���u�u�u�u�2�.��������F9��Y��D��4�
�:�&��+�(���Y����l�N��U���u�u�u�<��)�1���5����P��_�� ��`�%�g�i�w��(�������r/��h�����_�u�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}� ���&����	��h_�����3�
�e�
�d�}�JϮ�I����P��S/��B���
�<�n�u�w�}�W���YӃ��Z ���*���d�a�
�d�j�<�(���
����9��N�����u�u�u�u�w�}�W�������l ��h"����
�=�
� �`�h���E�Ƽ�9��D�����
�
�;�&�0�W�W���Y���F��D��]¡�%�3�
�f�`�-�W���	����@��AZ��\���=�;�_�u�w�}�W���Y���Z1��C1�����:�
�c�%�>�;�(��&����[��h^�����9�1��`�>����Y���F�N�����u�}�8�
�"�l�C؁�H����C9��Y�����a�|�!�0�w�}�W���Y���F������:�
�:�%�f���������l��R����� �&�4�0���(���
����F�N��U���0�&�3�}�#�-����J�ѓ�F�V�����
�#�
�|�w�5��ԜY���F�N��Uʼ�
�!��'��2�(���	����F9��1��G��u�
�
�;�4�1����J����@��=N��U���u�u�u�9�>�}�_���&���� R��G_��U���6�;�!�9�c�o�^Ϫ���ƹF�N��U���u�u��9��2�(���	����C��Q��Eߊ�f�u�h�%�g���������9��h��N���u�u�u�u�w�8����Qے��l ��]�*��h�4�
�:�$��ہ�P�Ƹ�V�N��U���u�u�u�u�>���������C9��h��*���b�`�%�g�k�}�(߁�����V��h_�����2�_�u�u�w�}�W������F�N��U���u�u�<�
�#���������l��h��B���%�g�i�u���/���!����k>��d��U���u�u�u�0�3�4�L���Y�����RNךU���u�u�u�u� �1�(���&����lW��G�����e�
�f�u�j��/���!����k>��o6�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u� �1�(���&����lW��G�����a�
�f�u�$�4�Ϯ�����F�=N��U���9�
�:�
�8�-�Fׁ�����lQ��h�*���<�;�%�:�w�}����
�μ�9��P�����e�<�
�<�{�-�B�������Z��h�����u�
�
�<�?�4����&����Z�G1��=����8�!�f�>����	�ӓ�Z��^��*ފ�;�&�2�u����������9��h��Yʥ�`��2��:�)�A���&������h&�����<�
�
�;�$�:�W���&������C1�����<�y�%�`��:�;����ߓ�]9��PB��*ߊ�<�=�<�<��m��������lS��^	�����
�d�<�
�>�q����1����Z��h_�����<�y�%�`��:�;�������Z��^	�����2��8�#�l�(���
���C9����9���!�d�
�;�$�:�W���&���� R��G_����<�
�1�
�d�m�W���
����W��Y����u�0�<�_�w�}�W����έ�l��h��*��c�u�=�;�w�}�W���Y����UF�C�����f�b�%�u�w�-��������lV����ߊu�u�u�u�w�}�W���.����u	��{��*���%�<�3�
�c��D���DӖ��l.��_"�����
�;�&�2�]�}�W���Y���V
��QN�����2�7�1�d�n�t����Y���F�N��U���u��9�
�8�����H˹��Z9��hY�*��u�h�%�`��:�;�������Z��^	�U���u�u�u�u�2�.��������F9��Y��D��4�
�:�&��+�(���Y����l�N��U���u�u�u�<��)�1���5����^��_�� ��g�%�g�i�w��(�������G9��h�����_�u�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}� ���&����	��h_�����3�
�a�
�d�}�JϮ�L����[*��^��F���
�<�n�u�w�}�W���YӃ��Z ���*���d�a�
�d�j�<�(���
����9��N�����u�u�u�u�w�}�W�������l ��h"����
�=�
� �`�o���E�Ƽ�9��P�����d�
�;�&�0�W�W���Y���F��D��]¡�%�3�
�f�`�-�W���	����@��AZ��\���=�;�_�u�w�}�W���Y���Z1��C1�����:�
�m�%�>�;�(��&����[��h[�����<�<�
�d�>����Y���F�N�����u�}�8�
�"�l�C؁�H����C9��Y������|�!�0�w�}�W���Y���F������:�
�:�%�f���������l��R������2��8�#�l�(���
����F�N��U���0�&�3�}�#�-����J�ѓ�F�V�����
�#�
�|�w�5��ԜY���F�N��Uʼ�
�!��'��2�(���	����F9��1��G��u�
�
�<�?�4����&����Z��N��U���u�u�0�&�1�u��������Q��N�����:�&�
�#��t�W������F�N��U���u�<�
�!��/�;���&�ޓ�[��B1�G���g�i�u�
��4��������Z��^	�U���u�u�u�u�2�.��������F9��Y��D��4�
�:�&��+�(���Y����l�N��U���u�u�u�<��)�1���5����^��_�� ��g�%�g�i�w��(�������G9��^ ����u�u�u�u�w�}��������^��B1�A݊�d�h�4�
�8�.�(���&���G��d��U���u�u�u�u�w�4�(���?����\	��V����� �b�g�%�e�a�W���&������C1�����<�n�u�u�w�}�W�������N��Z�� ��a�
�d�h�6�����&����O�C��U���u�u�u�u�w�}�WϷ�&����\��X��DҊ�=�
� �b�e�-�E��Y����{��{�����<�
�<�n�w�}�W���Y����_��F����� �d�a�
�f�`��������_��G�����u�u�u�u�w�}�W���Yӏ��_��X�����d�
�=�
�"�j�E���K���C9����9���!�a�<�
�>�f�W���Y���F��[��U���8�
� �d�c��F������]��[��F���!�0�u�u�w�}�W���Y�����[�����:�%�d�
�?����K����Z�G1��=����8�!�f�>����Y���F�N�����u�}�8�
�"�l�C؁�H����C9��Y�����g�|�!�0�w�}�W���Y���F������:�
�:�%�f���������l��R������2��8�#�o������ƹF�N��U���9�<�u�}�:����MĹ��[��G1�����9�a�d�|�#�8�W���Y���F�N��U���9�
�:�
�8�-�Fׁ�����lQ��h�U��%�`��2��0��������T]ǻN��U���u�u�9�0�]�}�W���Y���F�^9�����'��:�
�o�-����&����CU��S��-���������U�ԜY���F�N��ʼ�n�u�u�u�w�8����Y���F�N��"���
�:�
�:�'�l�(���&����T��\��H���������/���B���F���U���u�u�u�0�3�-����
��ƓF�C��"���
�:�
�:�'�o�(���&����_��\�����;�%�:�0�$�}�Z���Yӏ��_��X�����g�
�=�
�"�j�N���K����Z��G��U���'�6�&�}����������l��D��U���
�:��8�#�l��������lQ��X�����g�<�
�<�{�-�@�������G9��^ �����%�b��"�>�4�(ہ�����F�� 1�����<�
�
�;�$�:�W���&����Z��hX�����2�u�
�
�8�����N����@����*����8�!�m�>����	�ѓ�\��Z��L���
�<�y�%�`�� �������l��D��U���
�:��8�#�l�(���
���C9��{�����
�g�<�
�>�q����5����^��]�����2�u�
�
�8�����Hǹ��l��N��B���"�<�<�
�b�4�(���UӒ��l ��]�*��u�%�&�2�5�9�F��UӇ��@��U
��D��|�u�u�7�0�3�W���Y����UF��G1�����1�d�b�|�#�8�}���Y���F�^��]���
� �d�a��l�JϿ�&����G9��1�\ʡ�0�u�u�u�w�}�W���Y����d9��h(��*���%�g�
�=��(�@���	���F�� 1�����<�
�
�;�$�:�}���Y���F�R�����%�&�2�7�3�l�N�������9F�N��U���u�u�u��;���������9��^1��*��
�f�u�h�'�j�;�������S��Y1���ߊu�u�u�u�w�}����Y�θ�C9��h_�B���u�u�%�6�9�)����<����[��=N��U���u�u�u�u�w�
��������\��1�����
�b�
�f�w�`����5����^��Z�����2�_�u�u�w�}�W�������N��G1��*��b�%�u�u�'�>�����ғ�O��_�����u�u�u�u�w�}�W�������A9��X��E���<�3�
�b��n�W��	�ѓ�\��Z��Dي�;�&�2�_�w�}�W���Y�Ʃ�@��F�����
�f�b�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����G9��E1�����e�%�<�3��j�(��Y����lQ��X�����d�
�;�&�0�W�W���Y���F��D��]¡�%�3�
�f�`�-�W���	����@��AZ��\���=�;�_�u�w�}�W���Y���Z1��C1�����:�
�e�%�>�;�(��&����[��hY�����8�!�d�
�9�.��ԜY���F�N�����}�!�%�3��n�@���Y�ƭ�l��D��ފ�|�u�=�;�]�}�W���Y���F�^9�����'��:�
�g�-����&����CU��S��*݊�:��8�!�f��������F�N��Uʰ�&�3�}�!�'�;�(��N����F��h�����#�
�|�u�?�3�}���Y���F�N�����!��'��8��G�������Q��G]�I���
�
�:��:�)�N���&����9F�N��U���u�9�<�u��0�(���H����CW������!�9�a�m�~�)����Y���F�N��U����9�
�:��2���&����U�� W��F���h�%�b�� �4����&����Z��N��U���u�u�0�&�1�u��������Q��N�����:�&�
�#��t�W������F�N��U���u�<�
�!��/�;���&�֓�[��B1�L���g�i�u�
��2�;����ѓ�]9��PUךU���u�u�u�u�;�4�W�������lW�� 1��U���%�6�;�!�;�i�A�������9F�N��U���u�u�u��;���������9��^1��*��
�f�u�h�'�j�;�������9��h��N���u�u�u�u�w�8����Qے��l ��]�*��h�4�
�:�$��ہ�P�Ƹ�V�N��U���u�u�u�u�>���������C9��h��*���b�l�%�g�k�}�(؁�����Z��h�����_�u�u�u�w�}�W������G��Q��F���%�u�u�%�4�3����M�����YNךU���u�u�u�u�w�}� ���&����	��h\�����3�
�b�
�d�}�JϮ�N������C1�����<�n�u�u�w�}�W�������N��Z�� ��a�
�d�h�6�����&���� O�C��U���u�u�u�u�w�}�WϷ�&����\��X��Gڊ�=�
� �b�n�-�E��Y����	��^��*ي�;�&�2�_�w�}�W���Y�Ʃ�@��F�����
�f�b�%�w�}��������ER��G�����_�u�u�u�w�}�W���Y����G9��E1�����e�%�<�3��j�(��Y����lQ��X�����g�<�
�<�l�}�W���Y�����^��]���
� �d�a��l�JϿ�&����G9��1�\ʡ�0�u�u�u�w�}�W���Y����d9��h(��*���%�g�
�=��(�@���	���F�� 1�����<�
�
�;�$�:�}���Y���F�R��U���u�u�u�u�w�}�WϷ�&����\��X��Gڊ�=�
� �b�n�-�E��YѾ��k>��o6��-����n�u�u�w�}�W�������U]ǻN��U���9�0�_�u�w�}�W���Y����G9��E1�����e�%�<�3��j�(��Y���k>��o6��-�����w�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����f��V��4���
�%�#�1�>�����
������T��[���_�u�u�
��3��������l��A�����<�
�&�<�9�-����Y����V��G1�� ���4�0��
��-����Y����f��V��4���
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����0��
�
�'�+��������9F�N��U���u�
�
�;�4�1����I����E
��^ �����h�%�e� �$�<����&ù��l��d��U���u�0�&�u�w�}�W���Y����lV��Y������e�4�
�;��������C9��b ������
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��m�����ƭ�@�������{�x�_�u�w��(�������r/��h�����4�&�2�
�%�>�MϮ�������h;�����1��e�u����������lV��E��U���
�;�6�9�3��G���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e� �&�4�2��(߁�	����O��_�����u�u�u�u�w��(�������r/��h�����i�u�
�
�9�>����0����F�N�����u�u�u�u�w�}�WϮ�I����P��S/��E���
�<�u�h�'�m�"�������z9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�"�������z9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��F߁�	����l��D�����2�
�'�6�m�-����
ۖ��l3��T�����d�
�%�#�3�}�(߁�����V��h_�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l3��T�����d�
�%�#�3�t����Y���F�N��U���
�;�6�9�3��F߁�	����l��D��I���
�
�;�6�;�9�>��&����_��N��U���0�&�u�u�w�}�W���YӖ��l3��T�����d�
�%�#�3�4�(���Y����lV��Y������d�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��l�(���
����@��YN�����&�u�x�u�w�-�G���
����W'��^�����2�4�&�2��/���	����@��h^�����9�1��d�{�-�G���
����W'��^�����u�
�
�;�4�1����Hù��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�9�>����0����R��[
��U���;�_�u�u�w�}�W���&ù��@��R
��*���<�
�<�u�j�-�G���
����W'��^�U���u�u�0�&�w�}�W���Y�����h;�����1��d�
�9�.���Y����f��V��4���e�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l3��T�����d�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������lW��V�����;�&�2�4�$�:�(�������A	��D��*ڊ�;�6�9�1��l�(������C9��b ������
�d�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ڊ�;�6�9�1��l�(��������YNךU���u�u�u�u����������lW��V�����;�&�2�i�w��(�������r/��1��*���n�u�u�u�w�8����Y���F�N��*ڊ�;�6�9�1��l�(�������]9��PN�U���
�;�6�9�3��Fށ�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��3��������9��h��U���<�;�%�:�2�.�W��Y����lV��Y������d�
�;�$�:��������\������}�
�
�;�4�1����H����lV��Y������d�
�'�0�}�(߁�����V��h_�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��v'��D���
�9�|�u�?�3�}���Y���F�G1�� ���4�0��
�f�4�(���Y����lV��Y������d�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�;�6�;�9�>��&����Z�
N��E���&�4�0���l����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��l�(�������]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���g�4�
�9��3��������]9��X��U���6�&�}�
��3��������9��h��Yʥ�e� �&�4�2��(�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��3��������9��h��\���=�;�_�u�w�}�W���Y����f��V��4���g�4�
�9��3����E�Ƽ�9��D�����
�g�4�
�;�f�W���Y����_��=N��U���u�u�u�
��3��������9��h��*���&�2�i�u����������lW��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��F݁�����l��^	�����u�u�'�6�$�u�(߁�����V��h_�U���
�;�6�9�3��F݁����C9��b ������
�g�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����0��
�g�6�����Y����l�N��U���u�%�e� �$�<����&�ԓ�]9��PN�U���
�;�6�9�3��F��Y���F��[�����u�u�u�u�w��(�������r/��1��*���u�h�%�e��.����8����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��3�������� 9��h��*���&�2�4�&�0�}����
���l�N��E���&�4�0���n��������l��h�����%�:�u�u�%�>����&ù��@��R
��*���4�
�9�y�'�m�"�������z9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��@��R
��*���4�
�9�|�w�5��ԜY���F�N��E���&�4�0���n��������l��R����� �&�4�0���D���&����9F�N��U���0�_�u�u�w�}�W���&ù��@��R
��*���4�
�9�
�9�.���Y����f��V��4���f�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
�d�4�(���Y����T��E�����x�_�u�u����������lW��^ �����&�<�;�%�8�}�W�������C9��b ������
�f�u����������lW��G��Yʥ�e� �&�4�2��(�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e� �&�6�8�6���J����E
��N�����u�u�u�u�w�}����,����_��~1�*���&�2�i�u����������lW��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��D�����
�f�<�
�>�}�JϮ�I����P��S/��Dي�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��@��R
��*���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e��.����8����l��A�����<�
�&�<�9�-����Y����V��G1�� ���4�0��
�c�<�(���UӖ��l3��T�����d�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�� ���4�0��
�c�<�(���P�Ƹ�V�N��U���u�u�%�e��.����8����l��A�����<�u�h�%�g���������R��G1���ߊu�u�u�u�;�8�}���Y���F�G1�� ���4�0��
�c�<�(���&����Z�
N��E���&�4�0���i��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�e� �$�<����&�ғ�]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���a�<�
�<��.����	����	F��X��¥�e� �&�4�2��(��Y����f��V��4���a�%�0�y�'�m�"�������z9��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G���
����W'��Z�����1�|�!�0�w�}�W���Y�����h;�����1��d�
�9�.���Y����f��V��4���a�_�u�u�w�}����s���F�N����� �&�4�0���C���&����[��h^�����9�1��d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
�b�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I����P��S/��Dߊ�%�#�1�<��4�(�������A	��N�����&�%�e� �$�<����&�ӓ�C9��SB��*ڊ�;�6�9�1��l�(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�e� �$�<����&�ӓ�C9��SG�����u�u�u�u�w�}�WϮ�I����P��S/��Dߊ�%�#�1�<��4�W��	�֓�]��[��<��
�%�#�1�]�}�W���Y����l�N��U���u�%�e� �$�<����&�ӓ�C9��S1��*���u�h�%�e��.����8����l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����,����_��~1�*���&�2�4�&�0�}����
���l�N��E���&�4�0���h��������@��h����%�:�0�&�'�m�"�������z9��N��E���&�4�0���h����UӖ��l3��T�����d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lV��Y������d�
�%�!�9�^Ϫ���ƹF�N��U���
�
�;�6�;�9�>��&����Z�
N��E���&�4�0���h�}���Y���V
��d��U���u�u�u�%�g���������S��Y1����u�
�
�;�4�1����Hƹ��V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�e� �$�<����&¹��l��h�����4�&�2�u�%�>���T���F��1�����0��
�
�'�+����&����R��P �����o�%�:�0�$�-�G���
����W'��1��*���y�%�e� �$�<����&¹��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�m�"�������z9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��D�����
�
�%�#�3�4�(���Y����lV��Y������d�4�
�;�f�W���Y����_��=N��U���u�u�u�
��3��������l��A�����<�u�h�%�g���������9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��v'��*���&�2�4�&�0�}����
���l�N��E���&�4�0�����������Z��G��U���'�6�&�}����������lW�G1�� ���4�0��
��/����&ù��@��R
��*ۊ�%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�֓�]��[��<���4�
�9�|�w�5��ԜY���F�N��E���&�4�0����������C9��b ������
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�;�6�;�9�>�������TF���*���6�9�1��f�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���6�9�1��e�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I����P��S/��G���
�9�
�;�$�:��������\������}�
�
�;�4�1����K����E
����*���6�9�1��e�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�;�6�;�9�>�������WO�C��U���u�u�u�u�w�-�G���
����W'��1��*���
�;�&�2�k�}�(߁�����V��h\�����1�_�u�u�w�}����s���F�N����� �&�4�0���(�������]9��PN�U���
�;�6�9�3��E���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e��.����8����Z��^	�����;�%�:�0�$�}�Z���YӖ��l3��T�����g�<�
�<��.����	����	F��X��¥�e� �&�4�2��(��	�֓�]��[��<���%�0�y�%�g���������9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u����������lT��G1�����!�0�u�u�w�}�W���YӖ��l3��T�����g�<�
�<�w�`����,����_��~1����u�u�u�9�2�W�W���Y���F��1�����0��
�
�9�.���Y����f��V��4���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����f��V��4���
�%�#�1�>�����
������T��[���_�u�u�
��3��������l��A�����<�
�&�<�9�-����Y����V��G1�� ���4�0��
��-����Y����f��V��4���
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����0��
�
�'�+��������9F�N��U���u�
�
�;�4�1����J����E
��^ �����h�%�e� �$�<����&����l��d��U���u�0�&�u�w�}�W���Y����lV��Y������f�4�
�;��������C9��b ������
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�;�6�9�1��n�����ƭ�@�������{�x�_�u�w��(�������r/��h�����4�&�2�
�%�>�MϮ�������h;�����1��f�u����������lU��E��U���
�;�6�9�3��D���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e� �&�4�2��(܁�	����O��_�����u�u�u�u�w��(�������r/��h�����i�u�
�
�9�>����0����F�N�����u�u�u�u�w�}�WϮ�I����P��S/��F���
�<�u�h�'�m�"�������z9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�"�������z9��V�����;�&�2�4�$�:�W�������K��N����� �&�4�0���(�������]9��P1�����
�'�6�o�'�2����	�֓�]��[��<���4�
�9�y�'�m�"�������z9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�I����P��S/��A���
�9�|�u�?�3�}���Y���F�G1�� ���4�0��
��-��������TF���*���6�9�1��c�<�(���B���F����ߊu�u�u�u�w�}�(߁�����V��hZ�����1�<�
�<�w�`����,����_��~1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��D�����
�
�;�&�0�<����Y����V��C�U���%�e� �&�6�8�6���&����Z��D�����:�u�u�'�4�.�_���&����R
��v'��Yʥ�e� �&�4�2��(ہ����C9��b ������
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h;�����1��a�4��1�^������F�N��U���%�e� �&�6�8�6���&����Z�
N��E���&�4�0���f�W���Y����_��=N��U���u�u�u�
��3��������l��D��I���
�
�;�6�;�9�>���	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�;�6�;�9�>�������W9��h��U���<�;�%�:�2�.�W��Y����lV��Y������`�4�
�;���������Z��G��U���'�6�&�}����������lS��G1�����
�
�;�6�;�9�>�������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��3��������l��A��\ʡ�0�u�u�u�w�}�W���	�֓�]��[��<���4�
�9�
�9�.���Y����f��V��4���
�%�#�1�]�}�W���Y����l�N��U���u�%�e� �$�<����&ƹ��l��h�����i�u�
�
�9�>����0�ӓ�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�G���
����W'��1��*���u�&�<�;�'�2����Y��ƹF��h^�����9�1��`�>�����
����l��TN����0�&�%�e��.����8������h;�����1��`�%�2�q����,����_��~1�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R
��v'��*���#�1�|�!�2�}�W���Y���F��h^�����9�1��`�>�����DӖ��l3��T�����`�_�u�u�w�}����s���F�N����� �&�4�0���(���
���F��1�����0��
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�����0��
�
�'�+����&����R��P �����&�{�x�_�w�}�(߁�����V��hX�����1�<�
�<��.����	����	F��X��¥�e� �&�4�2��(ف�	����F��1�����0��
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N����� �&�4�0���(��������YNךU���u�u�u�u����������lP��G1�����
�<�u�h�'�m�"�������z9��V����u�u�u�u�2�.�W���Y���F���*���6�9�1��a�<�(���&����Z�
N��E���&�4�0�����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�;�4�1����O����@��V�����'�6�&�{�z�W�W���&ù��@��R
��*܊�;�&�2�4�$�:�(�������A	��D��*ڊ�;�6�9�1��k�W���&����R
��v'��*���2�u�
�
�9�>����0�Г�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�e��.����8����R��[
��U���;�_�u�u�w�}�W���&ù��@��R
��*܊�;�&�2�i�w��(�������r/��d��U���u�0�&�u�w�}�W���Y����lV��Y������c�<�
�>�}�JϮ�I����P��S/��C���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�I����P��S/��B���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�e� �$�<����&Ĺ��l��h�����4�&�2�
�%�>�MϮ�������h;�����1��b�4��1�[Ϯ�I����P��S/��B���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lV��Y������b�4�
�;�t�W������F�N��Uʥ�e� �&�4�2��(؁�	����l��D��I���
�
�;�6�;�9�>�������W]ǻN��U���9�0�_�u�w�}�W���Y����f��V��4���
�%�#�1�>�����DӖ��l3��T�����b�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�� ���4�0��
��3��������]F��X�����x�u�u�%�g���������9��h��*���<�;�%�:�w�}����
�μ�9��D�����
�y�%�e��.����8����C��N��E���&�4�0����������F��P��U���u�u�<�u��-��������Z��S��*ڊ�;�6�9�1��j�������G��d��U���u�u�u�%�g���������9��h��U��%�e� �&�6�8�6���B���F����ߊu�u�u�u�w�}�(߁�����V��hY�����2�i�u�
��3��������l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��3��������l��A�����<�u�&�<�9�-����
���9F���*���6�9�1��o�<�(���&����Z��D�����:�u�u�'�4�.�_���&����R
��v'��*���#�1�u�
��3��������l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(߁�����V��hV�����1�|�!�0�w�}�W���Y�����h;�����1��m�4��1�(���
���F��1�����0��
�
�'�+��ԜY���F��D��U���u�u�u�u�'�m�"�������z9��V�����;�&�2�i�w��(�������r/��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�֓�]��[��<���<�
�<�u�$�4�Ϯ�����F�=N��U���
�;�6�9�3��O���&����R��P �����o�%�:�0�$�-�G���
����W'��B��*ڊ�;�6�9�1��e����UӖ��l3��T�����m�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��D�����
�
�%�#�3�t����Y���F�N��U���
�;�6�9�3��O���&����[��h^�����9�1��m�]�}�W���Y����l�N��U���u�%�e� �$�<����&˹��l��R����� �&�4�0���(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C���� �&�4�0���(�������]9��PN�����u�'�6�&�y�p�}���Y����f��V��4���
�%�#�1�>�����
����l��TN����0�&�%�e��.����8����R��[
���� �&�4�0���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�e� �$�<����&ʹ��l��G�����_�u�u�u�w�}�W���&����R
��v'��*���#�1�<�
�>�}�JϮ�I����P��S/��L���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�;�6�;�9�>�������W9��h��U��%�e� �&�6�8�6���&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u����������l_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��b ������
�
�;�$�:��������\������}�
�
�;�4�1����@�Ƽ�9��D�����
�
�'�2�w��(�������r/��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G���
����W'��1��*���|�u�=�;�]�}�W���Y���C9��b ������
�
�;�$�:�K���&ù��@��R
��*��u�u�u�u�2�.�W���Y���F���*���6�9�1��n�4�(���Y����lV��Y������l�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W���	����f��V��9���!�<�=� �w�`����
����9��Q��C���%�b�_�u�w�p�W���I����P��S"�����2��!�4��1�W�������A	��D�X�ߊu�u�
�e��.����5����{��x�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���K����lW�R�����b�3�
�f�b�-�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g�1�0�F����Ƣ�GN��G1�����9�d�e�h�2�4����N����U��h�\���!�0�u�u�w�}�W���YӖ��9��D�����8�!�<�=�"��������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�e� �&�6�8�;�������|��V�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���d� �&�4�2���������R��[
�����2�4�&�2�w�/����W���F�G1�*���6�9�1�<�>�� �������W9��h��*���<�;�%�:�w�}����
�μ�W��Y�����<�<��"�9�<�(���UӖ��9��D�����8�!�:���-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�d�
�;�6�;�9����5����l��A��\ʡ�0�u�u�u�w�}�W���	����f��V��9���!�:��
�'�+����&����[��h_�� ���4�0��8�#�2�>���	����l�N��Uʰ�&�u�u�u�w�}�W���	����f��V��9���!�:��
�'�+����&����[��h_�� ���4�0��8�#�2�>���	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
�f���������Z��@'�����<�u�&�<�9�-����
���9F���D���&�4�0��:�)����&����Z��D�����:�u�u�'�4�.�_���H����P��S"�����"�;�u�
�f���������Z��@'�����y�%�d�
�9�>��������\��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�Fށ�����V��Z�����
�%�#�1�~�)����Y���F�N��*��� �&�4�0��0����0����l��R����
�;�6�9�3�4��������F�N�����u�u�u�u�w�}�WϮ�H¹��@��R
�����:��
�;�$�:�K���&�ד�]��[������"�;�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����1�����<�<�
�%�!�9�����ƭ�@�������{�x�_�u�w��E�������^��V�����;�&�2�4�$�:�(�������A	��D��*����0�'�<�>������Ƽ�T��[��9���!�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_��6���'�<�<�
�'�+��������9F�N��U���u�
�g��2�/����&����_��Y1����u�
�g��2�/����&����_��N��U���0�&�u�u�w�}�W���YӖ��9��R�����
�%�#�1�>�����DӖ��9��R�����
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h_��6���'�<�<�
�9�.�Ͽ�
����C��R��U���u�u�%�d��1��������]9��P1�����
�'�6�o�'�2����	����p
��E"�����%�d�
�9�6�����	������1�����<�<�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������1�����<�<�
�%�!�9�^Ϫ���ƹF�N��U���
�g��0�%�4��������Z�G1�*���4��8�!�]�}�W���Y����l�N��U���u�%�d�
�;�<�;�������@��S��*����0�'�<�>�����s���F�R ����_�u�u�;�w�/����B���F��\������8�!�'�6���������9��R��]��%�d�
�9�6���������TJ��C����x�|�_�u�w��B���
����W*��^�����u�h�%��$�1�(ف�&����^��G_����u�x�u�
�b���������Z��@!��*���#�1�4�&�0�}����
���l�N��Dߊ�;�6�9�1�>�4�;�������l��h�����%�:�u�u�%�>����	������D�����
��&�g�1�0�F�������]��Q��F���%�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��G���8�d�u�;�w�2�_ǿ�&����G9��1�Hʰ�<�6�;�b�1��D���	���F��R ��U���u�u�u�u�'�l�(���������C"��:���4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��h;�����1�<�<�� �(�(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l*��^�����0�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������_��V�����;�&�2�4�$�:�(�������A	��D��*ۊ�<�<�<�;�5�8�(������C9��{�����4�9�1�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ۊ�<�<�<�;�5�8�(��������YNךU���u�u�u�u����������_��V�����;�&�2�i�w��(�������R��S1��*���n�u�u�u�w�8����Y���F�N��*ۊ�<�<�<�;�5�8�(�������]9��PN�U���
�<�<�<�9�?����	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��4��������W9��h��U���<�;�%�:�2�.�W��Y����lW��^�����7�0�
�;�$�:��������\������}�
�
�<�>�4��������lW��^�����7�0�
�'�0�}�(ށ�����v��[�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����G��V�����
�9�|�u�?�3�}���Y���F�G1��9���!��4�9�3�4�(���Y����lW��^�����7�0�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�<�<�>�3����&����Z�
N��D���8�!��4�;�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�<�=�<�<����������@��V�����'�6�&�{�z�W�W���&ƹ��T��Z��E���
�9�
�;�$�:��������\������}�
�
�<�?�4����&����_�G1��=����8�!�e�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�<�=�<�>��(��������YNךU���u�u�u�u����������9��h��*���&�2�i�u����������9��h��N���u�u�u�0�$�}�W���Y���F��h[�����<�<�
�
�'�+����&����[��h[�����<�<�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�<�=�<�>��(���
����@��YN�����&�u�x�u�w�-�B�������Z��h�����4�&�2�
�%�>�MϮ�������h&�����<�
�y�%�b���������l��PB��*ߊ�<�=�<�<���������F��P��U���u�u�<�u��-��������Z��S��*ߊ�<�=�<�<����������[��=N��U���u�u�u�
��4��������Z��^	��Hʥ�`��2��:�)�G�ԜY���F��D��U���u�u�u�u�'�h�?���5����lV��Y1����u�
�
�<�?�4����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�`��2��0���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9����9���!�d�
�%�!�9��������@��h����%�:�0�&�'�h�?���5����lW��V�����%�`��2��0���&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�b���������9��h��\���=�;�_�u�w�}�W���Y����{��{����
�%�#�1�>�����DӖ��l.��_"�����e�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
�>�5����&�֓�C9��S1��*���u�h�%�`��:�;�������R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ځ�����^��^�����2�4�&�2�w�/����W���F�G1��=����8�!�d��3��������]9��X��U���6�&�}�
��4��������F��1�����8�!�d�
�%�:�W���&������C1�*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�L����[*��^��E���
�9�|�u�?�3�}���Y���F�G1��=����8�!�d��3����E�Ƽ�9��P�����d�n�u�u�w�}����Y���F�N��U���
�<�=�<�>��G���&����[��h[�����<�<�
�e�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h[�����<�<�
�d�6�����������^	�����0�&�u�x�w�}����1����Z��h_�����9�
�;�&�0�<����&����\��E�����
�
�<�=�>�4�(�������WJ��h[�����<�<�
�d�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�<�=�<�>��F���&����F��R ��U���u�u�u�u�'�h�?���5����lW��V�����;�&�2�i�w��(�������G9��h�����_�u�u�u�w�1��ԜY���F�N��@���2��8�!�f���������@��S��*ߊ�<�=�<�<��l��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�`��0�����H¹��l�������%�:�0�&�w�p�W���	�ӓ�Z��^��*���<�
�<�
�$�4��������C��R������2��8�#�l�[Ϯ�L����[*��^��D���0�y�%�`��:�;�������R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��4��������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�Z��^��*���<�
�<�u�j�-�B�������Z��UךU���u�u�9�0�]�}�W���Y���C9����9���!�d�
�;�$�:�K���&ƹ��T��Z��Dۊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ƹ��T��Z��D؊�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�>�5����&�ԓ�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����8�!�d�
�'�+����&ƹ��T��Z��D؊�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9����9���!�d�
�%�!�9�^Ϫ���ƹF�N��U���
�
�<�=�>�4�(�������W9��h��U��%�`��2��0���&����_��N��U���0�&�u�u�w�}�W���YӖ��l.��_"�����g�4�
�9��3����E�Ƽ�9��P�����d�
�%�#�3�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���=�<�<�
�e�4�(���Y����T��E�����x�_�u�u����������T��Y1�����&�2�
�'�4�g��������lS��^	�����
�g�u�
��4��������l��PB��*ߊ�<�=�<�<��o������ƹF��R	�����u�u�u�3��<�(���
����T��N������2��8�#�l�(��������YNךU���u�u�u�u����������T��Y1����u�
�
�<�?�4����K���F�N�����u�u�u�u�w�}����1����Z��h_�����<�u�h�%�b���������9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�b��������� 9��h��*���&�2�4�&�0�}����
���l�N��@���2��8�!�f���������@��V�����'�6�o�%�8�8�Ǯ�L����[*��^��F���
�9�y�%�b��������� 9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����1����Z��h_�����9�|�u�=�9�W�W���Y���F��1�����8�!�d�
�'�+����&����[��h[�����<�<�
�f�6����Y���F��[�����u�u�u�u�w��(�������G9��h�����<�
�<�u�j�-�B�������Z��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����{��{����
�;�&�2�6�.��������@H�d��Uʥ�`��2��:�)�F܁�����l��^	�����u�u�'�6�$�u�(ځ�����^��]�����2��8�#�l�(����Ƽ�9��P�����d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lS��^	�����
�f�4�
�;�t�W������F�N��Uʥ�`��2��:�)�F܁�����Z�G1��=����8�!�d�l�}�W���YӃ��VFǻN��U���u�u�
�
�>�5����&�Փ�]9��PN�U���
�<�=�<�>��D�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�<�=�<�>��C���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l.��_"�����a�4�
�9��3��������]9��X��U���6�&�}�
��4��������l��A��U���
�<�=�<�>��C���&����C��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�>�5����&�ғ�C9��SG�����u�u�u�u�w�}�WϮ�L����[*��^��A���
�9�
�;�$�:�K���&ƹ��T��Z��Dފ�%�#�1�_�w�}�W������F�N��U���%�`��2��0���&����_��Y1����u�
�
�<�?�4����M����E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h�?���5����lW��^ �����&�<�;�%�8�8����T�����h&�����<�
�a�<��4�(�������A	��N�����&�%�`��0�����H����lS��^	�����
�a�%�0�{�-�B�������Z��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ځ�����^��Z�����1�|�!�0�w�}�W���Y�����h&�����<�
�a�<��4�W��	�ӓ�Z��^��*��_�u�u�u�w�1��ԜY���F�N��@���2��8�!�f��������C9����9���!�d�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9����9���!�d�
�%�!�9�����ƭ�@�������{�x�_�u�w��(�������G9��h�����<�
�<�
�$�4��������C��R������2��8�#�l�(������C9����9���!�d�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��@���2��8�!�f���������[��=N��U���u�u�u�
��4��������l��A�����<�u�h�%�b���������9��h��N���u�u�u�0�$�}�W���Y���F��h[�����<�<�
�`�6���������Z�G1��=����8�!�d��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�<�=�>�4�(�������TF��D��U���6�&�{�x�]�}�W���&������C1�*���&�2�4�&�0�����CӖ��P����*���=�<�<�
�b�}�(ځ�����^��[�����u�
�
�<�?�4����L����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�`��0�����Hƹ��l��G�����_�u�u�u�w�}�W���&������C1�*���&�2�i�u����������S��N��U���0�&�u�u�w�}�W���YӖ��l.��_"�����`�<�
�<�w�`����1����Z��h_�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����1����Z��h_�����1�<�
�<�w�.����	����@�CךU���
�
�<�=�>�4�(ށ�	����l��D�����2�
�'�6�m�-����
ۖ��l.��_"�����
�%�#�1�w��(�������G9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�L����[*��^��*���#�1�|�!�2�}�W���Y���F��h[�����<�<�
�
�'�+����&����[��h[�����<�<�
�
�'�+��ԜY���F��D��U���u�u�u�u�'�h�?���5����lW��G1�����
�<�u�h�'�h�?���5����lW��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�L����[*��^��*���&�2�4�&�0�}����
���l�N��@���2��8�!�f�4�(���&����T��E��Oʥ�:�0�&�%�b���������F��1�����8�!�d�%�2�q����1����Z��h_�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����1����Z��h_�����1�|�!�0�w�}�W���Y�����h&�����<�
�
�;�$�:�K���&ƹ��T��Z��D�ߊu�u�u�u�;�8�}���Y���F�G1��=����8�!�d�>�����DӖ��l.��_"�����
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����{��{�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�`��:�;����ԓ�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����8�!�g�4��1�[Ϯ�L����[*��^��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��P�����g�4�
�9�~�}����s���F�N������2��8�#�o��������l��R������2��8�#�o������ƹF�N�����_�u�u�u�w�}�W���&������C1�����9�
�;�&�0�a�W���&������C1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��P�����g�<�
�<�w�.����	����@�CךU���
�
�<�=�>�4�(݁�����l��^	�����u�u�'�6�$�u�(ځ�����^��B��*ߊ�<�=�<�<������Y����{��{�����4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����{��{�����4�
�9�|�w�5��ԜY���F�N��@���2��8�!�e�4�(���Y����lS��^	�����
�n�u�u�w�}����Y���F�N��U���
�<�=�<�>��(���
���F��1�����8�!�g�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h&�����<�
�
�%�!�9�����ƭ�@�������{�x�_�u�w��(�������G9��V�����;�&�2�4�$�:�(�������A	��D��*ߊ�<�=�<�<�������Ƽ�9��P�����f�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h[�����<�<�
�
�'�+��������9F�N��U���u�
�
�<�?�4����&����_��Y1����u�
�
�<�?�4����&����_��N��U���0�&�u�u�w�}�W���YӖ��l.��_"�����
�%�#�1�>�����DӖ��l.��_"�����
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h[�����<�<�
�
�9�.�Ͽ�
����C��R��U���u�u�%�`��:�;����Փ�]9��P1�����
�'�6�o�'�2����	�ӓ�Z��^��*���%�`��2��0����	������h&�����<�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h&�����<�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�<�=�>�4�(܁�����Z�G1��=����8�!�f�]�}�W���Y����l�N��U���u�%�`��0�����J����@��S��*ߊ�<�=�<�<������s���F�R ����_�u�u�;�w�/����B��ƹF�N��@���2��8�!�c�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L����[*��^��*���#�1�<�
�>���������PF��G�����%�`��2��0��������WJ��h[�����<�<�
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N������2��8�#�i�������G��d��U���u�u�u�%�b���������l��A�����<�u�h�%�b���������l��A�����u�u�u�9�2�W�W���Y���F��1�����8�!�a�4��1�(���
���F��1�����8�!�a�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����2��8�#�i�����ƭ�@�������{�x�_�u�w��(�������G9��^ �����&�<�;�%�8�}�W�������C9����9���!�a�u�
��4��������C��N��@���2��8�!�c�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��@���2��8�!�c�<�(���P�Ƹ�V�N��U���u�u�%�`��:�;����ғ�]9��PN�U���
�<�=�<�>��L���Y�����RNךU���u�u�u�u����������9��h��U��%�`��2��0����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�<�=�>�4�(ځ�	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��P�����`�4�
�9��3��������]9��X��U���6�&�}�
��4��������R��[
�����2��8�#�h��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�<�?�4����&����_����ߊu�u�u�u�w�}�(ځ�����^��1��*���
�;�&�2�k�}�(ځ�����^��1��*���n�u�u�u�w�8����Y���F�N��*ߊ�<�=�<�<����������@��S��*ߊ�<�=�<�<����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�<�?�4����&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L����[*��^��*���&�2�4�&�0�����CӖ��P����*���=�<�<�
�{�-�B�������Z��h�����
�
�<�=�>�4�(ځ�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�<�=�>�4�(ځ�	����O��_�����u�u�u�u�w��(�������G9��^ �����h�%�`��0�����L���F�N�����u�u�u�u�w�}����1����Z��h[�����2�i�u�
��4��������C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`��:�;����Г�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h[�����<�<�
�
�'�+����&����R��P �����o�%�:�0�$�-�B�������Z��h�����u�
�
�<�?�4����&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�b���������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�Z��^��*܊�%�#�1�<��4�W��	�ӓ�Z��^��*܊�%�#�1�_�w�}�W������F�N��U���%�`��2��0��������W9��h��U��%�`��2��0��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�b���������l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��P�����c�<�
�<��.����	����	F��X��¥�`��2��:�)�A���&ƹ��T��Z��C���0�y�%�`��:�;����Г�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�`��:�;����Г�C9��SG�����u�u�u�u�w�}�WϮ�L����[*��^��*���&�2�i�u����������]ǻN��U���9�0�_�u�w�}�W���Y����{��{�����<�
�<�u�j�-�B�������Z��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������G9��V�����;�&�2�4�$�:�W�������K��N������2��8�#�j��������l��h�����%�:�u�u�%�>����&ƹ��T��Z��B���
�9�y�%�b���������l��A�����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ځ�����^�� 1��*���|�u�=�;�]�}�W���Y���C9����9���!�b�4�
�;��������C9����9���!�b�4�
�;�f�W���Y����_��=N��U���u�u�u�
��4��������R��[
�����2�i�u�
��4��������R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ځ�����^�� 1��*���u�&�<�;�'�2����Y��ƹF��h[�����<�<�
�
�9�.����
����C��T�����&�}�
�
�>�5����&����lS��^	�����
�
�'�2�w��(�������G9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(�������G9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��P�����b�<�
�<�w�`����1����Z��hY�U���u�u�0�&�w�}�W���Y�����h&�����<�
�
�;�$�:�K���&ƹ��T��Z��B���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�L����[*��^��*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�<�?�4����&����_��Y1�����&�2�
�'�4�g��������lS��^	�����
�
�%�#�3�}�(ځ�����^��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ӓ�Z��^��*Ҋ�%�#�1�|�#�8�W���Y���F���*���=�<�<�
��-��������TF���*���=�<�<�
��-����s���F�R��U���u�u�u�u�w�-�B�������Z��h�����<�
�<�u�j�-�B�������Z��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�Z��^��*Ҋ�;�&�2�4�$�:�W�������K��N������2��8�#�e��������@��h����%�:�0�&�'�h�?���5����l^�G1��=����8�!�m�'�8�[Ϯ�L����[*��^��*���#�1�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�L����[*��^��*���#�1�|�!�2�}�W���Y���F��h[�����<�<�
�
�9�.���Y����{��{����_�u�u�u�w�1��ԜY���F�N��@���2��8�!�o�4�(���Y����lS��^	�����
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��P�����l�4�
�9��3��������]F��X�����x�u�u�%�b���������l��A�����<�
�&�<�9�-����Y����V��G1��=����8�!�l�6����	�ӓ�Z��^��*ӊ�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9����9���!�l�4�
�;�t�W������F�N��Uʥ�`��2��:�)�N���&����Z��^	��Hʥ�`��2��:�)�N���&����9F�N��U���0�_�u�u�w�}�W���&ƹ��T��Z��L���
�9�
�;�$�:�K���&ƹ��T��Z��L���
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9����9���!�l�<�
�>�}����Ӗ��P��N����u�
�
�<�?�4����&����Z��D�����:�u�u�'�4�.�_���&������C1�U���
�<�=�<�>��(����Ƽ�9��P�����l�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��P�����l�4�
�9�~�}����s���F�N������2��8�#�d���������h&�����<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�<�=�>�4�(ց�����Z�G1��=����8�!�l�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY�����8�!�e�4��1�(���
����@��YN�����&�u�x�u�w�-�@�������G9��V�����;�&�2�4�$�:�(�������A	��D��*݊�:��8�!�g�<�(���UӖ��l*��{�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h"��9���!�e�4�
�;�t�W������F�N��Uʥ�b��"�<�>��(�������]9��PN�U���
�:��8�#�m������ƹF�N�����_�u�u�u�w�}�W���&����Z��h^�����1�<�
�<�w�`����5����^��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����	��^��*ڊ�;�&�2�4�$�:�W�������K��N������"�<�<����������Z��G��U���'�6�&�}����������F�� 1�����<�
�
�'�0�}�(؁�����Z��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@�������G9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��@"�����
�;�&�2�k�}�(؁�����Z��d��U���u�0�&�u�w�}�W���Y����lQ��X�����e�<�
�<�w�`����5����^��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@�������G9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�:��8�#�l�(�������]9��P1�����
�'�6�o�'�2����	�ѓ�\��Z��Dڊ�%�#�1�u����������9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����5����^��^�����1�|�!�0�w�}�W���Y�����h"��9���!�d�
�%�!�9���������h"��9���!�d�
�%�!�9�}���Y���V
��d��U���u�u�u�%�`�� �������l��A�����<�u�h�%�`�� �������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����5����^��^�����2�4�&�2�w�/����W���F�G1��9���<�<�
�e�>�����
����l��TN����0�&�%�b��*����&���C9��{�����
�e�%�0�{�-�@�������G9��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@�������G9��h�����|�!�0�u�w�}�W���Y����lQ��X�����d�
�;�&�0�a�W���&����Z��h_����u�u�u�9�2�W�W���Y���F�� 1�����<�
�e�<��4�W��	�ѓ�\��Z��Dڊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&Ĺ��D*��^��D���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�b�� �4����H����E
��^ �����&�<�;�%�8�}�W�������C9��{�����
�d�4�
�;�q����5����^��_�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����	��^��*���4�
�9�|�w�5��ԜY���F�N��B���"�<�<�
�f�<�(���&����Z�
N��B���"�<�<�
�f�<�(���B���F����ߊu�u�u�u�w�}�(؁�����Z��1��*���
�;�&�2�k�}�(؁�����Z��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����	��^��*���<�
�<�u�$�4�Ϯ�����F�=N��U���
�:��8�#�l�(���
����@��Y1�����u�'�6�&���(���5����lW����*����8�!�d��/����&Ĺ��D*��^��D���
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��D*��^��D���
�9�|�u�?�3�}���Y���F�G1��9���<�<�
�d�>�����DӖ��l*��{����n�u�u�u�w�8����Y���F�N��*݊�:��8�!�f��������C9��{�����
�d�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lQ��X�����d�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������9��h��*���&�2�4�&�0�����CӖ��P����*����8�!�d��-����Y����	��^��*���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h"��9���!�d�
�%�!�9�^Ϫ���ƹF�N��U���
�
�:��:�)�F݁�	����l��D��I���
�
�:��:�)�F݁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�\��Z��D؊�%�#�1�<��4�W��	�ѓ�\��Z��D؊�%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h"��9���!�d�
�;�$�:�����Ƽ�\��D@��X���u�%�b�� �4����K����@��V�����'�6�o�%�8�8�Ǯ�N������C1�Yʥ�b��"�<�>��E�������lQ��X�����d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lQ��X�����d�
�%�#�3�t����Y���F�N��U���
�:��8�#�l�(���
���F�� 1�����<�
�g�_�w�}�W������F�N��U���%�b��"�>�4�(�������TF���*����8�!�d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��9���<�<�
�f�6�����������^	�����0�&�u�x�w�}����5����^��]�����1�<�
�<��.����	����	F��X��¥�b��"�<�>��D���&������h"��9���!�d�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��B���"�<�<�
�d�<�(���P�Ƹ�V�N��U���u�u�%�b��*����&�Փ�C9��S1��*���u�h�%�b��*����&�Փ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��{�����
�f�4�
�;��������C9��{�����
�f�4�
�;�����s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���"�<�<�
�d�4�(���Y����T��E�����x�_�u�u���������� 9��h��*���<�;�%�:�w�}����
�μ�9��@"�����f�u�
�
�8�����H����V�G1��9���<�<�
�f�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��9���<�<�
�f�6�����Y����l�N��U���u�%�b�� �4����J����@��S��*݊�:��8�!�f�f�W���Y����_��=N��U���u�u�u�
��2�;�������Z��^	��Hʥ�b��"�<�>��D�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�:��8�#�l�(�������]9��PN�����u�'�6�&�y�p�}���Y����	��^��*���4�
�9�
�9�.����
����C��T�����&�}�
�
�8�����Hǹ��l��N��B���"�<�<�
�c�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�:��:�)�Fہ�	����O��_�����u�u�u�u�w��(���5����lW��V�����;�&�2�i�w��(���5����lW��V����u�u�u�u�2�.�W���Y���F���*����8�!�d��-��������TF���*����8�!�d��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�:��:�)�Fہ�������^	�����0�&�u�x�w�}����5����^��Z�����2�4�&�2��/���	����@��hY�����8�!�d�y�'�j�;�������R��E��U���
�:��8�#�l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�:��8�#�l�(��������YNךU���u�u�u�u����������9��h��U��%�b��"�>�4�(��s���F�R��U���u�u�u�u�w�-�@�������G9��h�����i�u�
�
�8�����Hǹ��V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�b�� �4����L����E
��^ �����&�<�;�%�8�8����T�����h"��9���!�d�
�%�!�9��������@��h����%�:�0�&�'�j�;�������S��G1�����
�
�:��:�)�Fځ�	����l��PGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�b��*����&�ӓ�C9��SG�����u�u�u�u�w�}�WϮ�N������C1�*���#�1�<�
�>�}�JϮ�N������C1�*���#�1�_�u�w�}�W������F�N��Uʥ�b��"�<�>��B���&����Z��^	��Hʥ�b��"�<�>��B���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b��*����&�ӓ�]9��PN�����u�'�6�&�y�p�}���Y����	��^��*���<�
�<�
�$�4��������C��R������"�<�<��h�W���&����Z��h_�����y�%�b�� �4����L����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�b�� �4����L����E
��N�����u�u�u�u�w�}����5����^��[�����2�i�u�
��2�;�������9F�N��U���0�_�u�u�w�}�W���&Ĺ��D*��^��@���
�<�u�h�'�j�;�������S��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u����������l��A�����<�u�&�<�9�-����
���9F���*����8�!�d�6���������l��^	�����u�u�'�6�$�u�(؁�����Z��h�����u�
�
�:��0��������W9��R	��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��2�;����ד�C9��SG�����u�u�u�u�w�}�WϮ�N������C1�����9�
�;�&�0�a�W���&����Z��h_�����1�_�u�u�w�}����s���F�N������"�<�<����������@��S��*݊�:��8�!�f�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b��"�>�4�(ށ�������^	�����0�&�u�x�w�}����5����^��1��*���
�&�<�;�'�2�W�������@N�� 1�����<�
�y�%�`�� �������C��N��B���"�<�<�
��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*����8�!�d�6�����Y����l�N��U���u�%�b�� �4����&����Z�
N��B���"�<�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�8�����H����@��S��*݊�:��8�!�f�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*����8�!�g�6�����������^	�����0�&�u�x�w�}����5����^��1��*���
�;�&�2�6�.���������T��]���
�:��8�#�o��������lQ��X�����g�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY�����8�!�g�4��1�^������F�N��U���%�b��"�>�4�(݁�	����l��D��I���
�
�:��:�)�E���&����9F�N��U���0�_�u�u�w�}�W���&Ĺ��D*��^��*���#�1�<�
�>�}�JϮ�N������C1�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��@"�����
�;�&�2�6�.��������@H�d��Uʥ�b��"�<�>��(���
����@��Y1�����u�'�6�&���(���5����lT�G1��9���<�<�
�
�%�:�W���&����Z��h\�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����5����^��1��*���|�u�=�;�]�}�W���Y���C9��{�����
�
�;�&�0�a�W���&����Z��h\�U���u�u�0�&�w�}�W���Y�����h"��9���!�g�<�
�>�}�JϮ�N������C1�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����5����^��1��*���
�;�&�2�6�.��������@H�d��Uʥ�b��"�<�>��(�������]9��P1�����
�'�6�o�'�2����	�ѓ�\��Z��F���
�9�y�%�`�� �������R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�@�������G9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��@"�����
�%�#�1�>�����DӖ��l*��{�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�:��0��������W9��h��U��%�b��"�>�4�(܁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��2�;����Փ�]9��PN�����u�'�6�&�y�p�}���Y����	��^��*ي�;�&�2�4�$�:�(�������A	��D��*݊�:��8�!�d�}�(؁�����Z��h�����
�
�:��:�)�D���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b��"�<�>��(��������YNךU���u�u�u�u����������l��D��I���
�
�:��:�)�D�ԜY���F��D��U���u�u�u�u�'�j�;������� 9��h��U��%�b��"�>�4�(܁�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b��"�<�>��(�������]9��PN�����u�'�6�&�y�p�}���Y����	��^��*ފ�%�#�1�<��4�(�������A	��N�����&�%�b�� �4����&����_�G1��9���<�<�
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N������"�<�<����������[��=N��U���u�u�u�
��2�;����ғ�C9��S1��*���u�h�%�b��*����&ǹ��l��d��U���u�0�&�u�w�}�W���Y����lQ��X�����a�4�
�9��3����E�Ƽ�9��@"�����
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY�����8�!�a�<��4�W�������A	��D�X�ߊu�u�
�
�8�����M����@��V�����'�6�o�%�8�8�Ǯ�N������C1�U���
�:��8�#�i����UӖ��l*��{�����4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����	��^��*ފ�%�#�1�|�#�8�W���Y���F���*����8�!�a�>�����DӖ��l*��{����_�u�u�u�w�1��ԜY���F�N��B���"�<�<�
��3����E�Ƽ�9��@"�����
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����	��^��*ߊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�8�����L����E
��^ �����&�<�;�%�8�}�W�������C9��{�����
�
�%�#�3�}�(؁�����Z��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��D*��^��*���#�1�|�!�2�}�W���Y���F��hY�����8�!�`�4��1�(���
���F�� 1�����<�
�
�%�!�9�}���Y���V
��d��U���u�u�u�%�`�� �������R��[
�����2�i�u�
��2�;����ӓ�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@�������G9��^ �����&�<�;�%�8�8����T�����h"��9���!�`�<�
�>���������PF��G�����%�b��"�>�4�(��	�ѓ�\��Z��@���0�y�%�b��*����&ƹ��l��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�
�
�8�����L����E
��N�����u�u�u�u�w�}����5����^��1��*���u�h�%�b��*����&��ƹF�N�����_�u�u�u�w�}�W���&����Z��h[�����2�i�u�
��2�;����ӓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�8�����O����E
��^ �����&�<�;�%�8�8����T�����h"��9���!�c�4�
�;���������Z��G��U���'�6�&�}����������l��A��U���
�:��8�#�k��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�:��0��������WO�C��U���u�u�u�u�w�-�@�������G9��V�����;�&�2�i�w��(���5����lP��G1���ߊu�u�u�u�;�8�}���Y���F�G1��9���<�<�
�
�'�+����&����[��hY�����8�!�c�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����"�<�<������Ӈ��Z��G�����u�x�u�u�'�j�;�������9��h��*���<�;�%�:�w�}����
�μ�9��@"�����y�%�b�� �4����&����F�� 1�����<�
�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h"��9���!�c�4�
�;�t�W������F�N��Uʥ�b��"�<�>��(���
���F�� 1�����<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�:��:�)�A���&����[��hY�����8�!�c�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h"��9���!�b�4�
�;�����Ӈ��Z��G�����u�x�u�u�'�j�;�������9��h��*���&�2�4�&�0�����CӖ��P����*����8�!�b�6����	�ѓ�\��Z��B���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lQ��X�����b�4�
�9�~�}����s���F�N������"�<�<����������@��S��*݊�:��8�!�`�<�(���B���F����ߊu�u�u�u�w�}�(؁�����Z��h�����<�
�<�u�j�-�@�������G9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&Ĺ��D*��^��*���&�2�4�&�0�}����
���l�N��B���"�<�<�
��3��������]9��X��U���6�&�}�
��2�;������C9��{�����
�
�'�2�w��(���5����lQ��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�j�;�������9��h��\���=�;�_�u�w�}�W���Y����	��^��*݊�;�&�2�i�w��(���5����lQ��N��U���0�&�u�u�w�}�W���YӖ��l*��{�����<�
�<�u�j�-�@�������G9��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�;�������9��h��*���&�2�4�&�0�}����
���l�N��B���"�<�<�
��-��������T9��D��*���6�o�%�:�2�.����5����^��1��*���y�%�b�� �4����&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`�� �������R��[
��U���;�_�u�u�w�}�W���&Ĺ��D*��^��*���#�1�<�
�>�}�JϮ�N������C1�����9�n�u�u�w�}����Y���F�N��U���
�:��8�#�e��������l��R������"�<�<����������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�:��0��������TF��D��U���6�&�{�x�]�}�W���&����Z��hV�����2�4�&�2��/���	����@��hY�����8�!�m�u����������l��PB��*݊�:��8�!�o�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��B���"�<�<�
��-����PӒ��]FǻN��U���u�u�
�
�8�����A����@��S��*݊�:��8�!�o�W�W���Y�Ʃ�@�N��U���u�u�%�b��*����&˹��l��R������"�<�<������s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���"�<�<�
��-��������TF��D��U���6�&�{�x�]�}�W���&����Z��hW�����1�<�
�<��.����	����	F��X��¥�b��"�<�>��(������C9��{�����
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��9���<�<�
�
�'�+��������9F�N��U���u�
�
�:��0��������W9��h��U��%�b��"�>�4�(ց�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�\��Z��L���
�9�
�;�$�:�K���&Ĺ��D*��^��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lQ��X�����l�<�
�<�w�.����	����@�CךU���
�
�:��:�)�N���&����R��P �����o�%�:�0�$�-�@�������G9����*����8�!�l�'�8�[Ϯ�N������C1�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����Z��hW�����1�|�!�0�w�}�W���Y�����h"��9���!�l�<�
�>�}�JϮ�N������C1����u�u�u�9�2�W�W���Y���F�� 1�����<�
�
�;�$�:�K���&Ĺ��D*��^��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w��(�������P��R��R��"�0�u�!�'�.����N�ѓ�F�V�����
�#�c�e�w�1����^��ƹF�N��M���8�!�0�6�2�����Ӈ��Z��G�����u�x�u�u�'�e�;�������[��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�E������V��T��B���
�f�`�%�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������C9��Y�����e�h�0�<�4�3�@���&����l��G�����u�u�u�u�w�}�WϮ�A����Z��V�����
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��Z�����0�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�"�������Z����<���%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�9�>��������Z��Y1��*���
�;�&�2�6�.���������T��]���
�;�6�9�3�4��������R��[
���� �&�4�0��0��������C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���������C&�����4�
�9�|�w�5��ԜY���F�N��L���&�4�0��:�)��������E
��^ �����h�%�l� �$�<��������T��h�����_�u�u�u�w�1��ԜY���F�N��L���&�4�0��:�)��������E
��^ �����h�%�l� �$�<��������T��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�]��[������2��
�9�.�Ͽ�
����C��R��U���u�u�%�l��.����5����{��~ �����2�4�&�2��/���	����@��hW�����9�1�<�<��:�>��	�ߓ�]��[������2��
�%�:�W���&����R
��{�����=�;�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��b ������8�!�<�?�3�������G��d��U���u�u�u�%�n���������Z��P��*���&�2�i�u����������^��^	���ߊu�u�u�u�;�8�}���Y���F�G1�� ���4�0��8�#�4��������TF���*���6�9�1�<�>�����&����l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����&�9�
�
��(�F��&����[�F��]���}�}�}�4�%�1�(���&����lT��[��@���
�l�u�u�%���������C9��h_��Dފ� �g�c�u�w�/�(���?����\	��Y��@��
� �g�g�w�}��������l*��G1�*���d�
� �g�o�}�W���&����\��X��G݊�`�d�
� �e�i�W�������l ��h"����
�`�d�
�"�o�G���Y����_��X�����g�
�`�l�1��A���_Ӈ��l
��q��9���
�b�d�
��(�E��Y�ƭ�A9��h(��*���%�g�
�`�`�;�(��P����A��C1�����:�
�b�d�����M���R��[�����:�%�g�
�b�h����L�����h��3����:�
�b�f����I���R��[�����:�%�g�
�b�l����J�����h��3����:�
�b�f��(���K���F��E1��*���
�:�%�g��h�D���&����@��E�����'��:�
�`�l�(ہ�����]ǻN��*��� �!�c�&�1��A���	���F�F��]���}�}�}�'��)�1���5����_��1�*���f�a�s�4�%�1�(���&����lT��[��A���
�`�|�s�6�/��������\��1�*���3�
�a�|�q�<����&����	��h\��Dߊ�g�3�
�a�~�{��������A9��X��L��
�d�3�
�d�t�QϿ�����u	��{��*���d�
�e�3��n�^�������G9��E1�����l�d�
�
�"�n�G���Y����_��X�����g�
�`�m�1��E���_Ӈ��l
��q��9���
�l�d�
��(�D��Y�ƭ�A9��h(��*���%�g�
�`�a�;�(��P����A��C1�����:�
�l�d�����M���R��[�����:�%�g�
�b�i����H�����h��3����:�
�l�f��(���J���F��E1��*���
�:�%�g��h�E���&����@��E�����'��:�
�n�l�(ށ�����F�V�����:�
�:�%�e��B���&����l�N�����
�f�b�%�w�`��������l*��G1�����c�d�a�x�f�9� ���Y����F�C�����
�b�b�%�w�`�_�������lP��h��D��
�d�u�'�'�����&ƹ��U��Z����n�u�u� ���2�������l ��^�*��i�u�u�u�w�}��������_��h^�����}�:�9�-�����&����P��G\��\��r�r�u�9�2�W�W���Y�Ƽ�W��Y�����<�<��"�9�4�(���B������V�