-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǑ[�������n� �2��2�������T��_�[���n� �0���s�"���0����wH��[Uװ���!�u�g��n�d����������h��A���d�<�_�0�2�4�W�ԜY�ƅ�F�N��U���o�;�0�0�w�`�G�ԜY�Ƃ�~9��v)��U���o�;�0�0�w�`�F�ԜY�ƨ�]W��~*��U���u�u�<�!�0�/�M���K���F��Y\��<���u�u�u�u�>�)����C����l�N��ي���u�u�w�}�������F��d��Uʱ�;�
���w�}�W�������V�
N�N���u�1�;�
��	�W���Y����]��R��H��n�u�u�1�9��>���Y���F��Y�����h�f�n�u�w�9�؁�0����F�N�����0�u�h�f�l�}�WϺ�˹��w2��N��U���;�0�0�u�j�n�L���Yӂ��
9��s:��U���u�o�;�0�2�}�J��B�����^��<���u�u�u�u�>�)����C����l�N��������u�w�}�M�������	[�UךU���<�d�
���}�W���Yɏ��V��T��F��u�u�1�;�d�
�3���Y���\��C����u�g�_�u�w�4�Fہ�0����F�N�����0�u�h�f�l�}�WϺ��ӓ�z"��N��U���<�!�2�'�m�}�E�ԜY�ƨ�]W��`'��=���u�u�o�;�2�8�W��J��ƹF��^ �*����u�u�u�w�4������� T��N�����
���u�w�}�W�������AF��]�N��'�u�_�u�w�4�F���C���@��[�����6�:�}�u�8�3���B�����N��O���u�!�
�:�>���������\��XN�N���u�1�;�u�w�4�Wϭ�����Z��R����1�"�!�u�~�W�W������\��N�����2�6�#�6�8�u�W������]ǻN�����u�o�;�u�#�����&����\�
�����e�n�u�u�3�3�W�������G��X	��*���!�'�e�1� �)�W���s���W��N�����&�1�9�2�4�+����Q�ƨ�D��^����u�<�m�u�m�3�W���&����P9��T��]���:�;�:�e�l�}�WϺ����	����*���<�
�0�!�%�m��������l�N����u�o�;�u�#�����&����\�
�����e�n�u�u�3�3�F���C���@��[�����6�:�}�u�8�3���B�����\��Uм�u�&�1�9�0�>��������W	��C��\�ߊu�u�<�d�w�}����
����\��h�����e�1�"�!�w�t�}���Y����F���U���
�:�<�
�2�)�������\F��d��Uʱ�;�`�u�o�9�}��������E��X��U���;�:�e�n�w�}����O���Z�D�����6�#�6�:��}�������9F�
��D���u�<�u�&�3�1��������AN��S�����|�_�u�u�8�)�W���C����@��[�����6�:�}�u�8�3���P���WF��C��N���'�=�!�6�"�8�����ơ�q ��vW��*ڊ� �
�c�:��8�C���Hӏ��F�C�� ���<�!�'�4�w�4����s���@��V�����u�o�&�1�;�:�������� F��@ ��U���_�u�u�x�;�+���
����_ǻN�����9�8�-�d�g�}�W�������T��A�����u�:�;�:�g�f�W���
����_F��O1��D���u�u�!�
�8�4�(��������Y��E��u�u�&�2�6�}����&���\��C
�����
�0�!�'�g�9� ���Y����F�D����� �
�
�u�w�g��������l��C��Eʱ�"�!�u�|�]�}�W�������F��hZ��U��&�1�9�2�4�+����Q�ƨ�D��^����u�<�;�9�:�%�F��Y����@��[�����6�:�}�u�8�3���B�����Y�����d�c�u�u�w�)�(�������P��^�����:�e�n�u�w�.����Y����9��N��U���
�:�<�
�2�)�������\F��d��U���u�0�0�u�w�4����s���@��V�� ���
�u�u�o�$�9��������G	��N�����u�|�_�u�w�4��������lW�N����9�2�6�#�4�2�_�������V�=N��U���;�9�8�-�e�o�W���Y����_	��T1�����}�u�:�;�8�m�L���Yӕ��]��Z��G��u�u�u�!��2��������V��X����n�u�u�x�w�8����Y����R
��N�����4�u� �
��}�W��
����\��h�����e�1�"�!�w�t�}���Y����R
��B��*���u�o�&�1�;�:��������F��@ ��U���_�u�u�x�;�+���
����_ǻN�����9�8�-�a�g�}�W�������T��A�����u�:�;�:�g�f�������_F�
��D��_�x��;�%�)�W�������_	��Td�����e�i�u�<�f�*��������[�I�����1�;�n�8�/�l�F��Y������YN����u�u�e�u�;�8����B����lW��R�����u�=�;�&�;�m�W���I�Ʃ�@��^ ����
�
�u�h�3�3�W���ӕ��V�
N��Rʰ�&�u�<�m�]�(�(ށ�Y����Z��@��U���}�|�h�r�p�8��������9��h_��U��1�;�d�"�2�}����P���A��[�����g�_� �
��}�JϺ�����[��D��E���u�e�u�9�2�9���s����9��S����u�=�;�&�;�m�W���I�Ʃ�@��^ �N�߇x��;�'�#�}����Y�Ơ�T��Z��G��i�u� �
��}����
���F�^�����u� �
�
�l�0����H���^��1����u�0�}�|�j�z�Pϻ�
�ơ�K9��U�� ���
�u�h�8�/�l�Cϩ��ƿ�_N��S��E���9�0�8�-�f�h�}���&����[��B��*���=�;�&�9�f�}�W��Y������h_��N�߇x��;�'�#�}����Y�Ơ�T��Z��F��i�u� �
��}����
���F�^�����u� �
�
�l�0����H���^��1����u�0�}�|�j�z�Pϻ�
�ơ�K9��UװX���0�0�4�0�;�+�������9��hZ��U��8�-�f�e� �8�W���Q���A����ʸ�-�f�d�_�z�}����ӊ��Z��X��I��� �
�
�n�]�3�W�������G��d