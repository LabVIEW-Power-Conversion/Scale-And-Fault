-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��l����}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���_�u�u�
����������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�Ƽ�9��V�����u������4�ԜY�Ƽ�9��N��U���
���
��	�%���Lӂ��]��G�U���%�e�g�4��1�W���7ӵ��l*��~-�U���%�e�f�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I�Փ�C9��SN�<����
���l�}�WϮ�I���/��d:��9�������w�l�W������]ǻN��*ڊ�
�%�#�1�m��W���&����p]ǻN��*ڊ�u�u�����0���/����aF�N�����u�|�_�u�w��(ځ�	����\��yN��1�����_�u�w��(���Y����g"��x)��*�����}�`�3�*����P���F��1�����9�u�u����;���:���F��1�Oʜ�u��
����2���+������Y��E��u�u�%�e�`�<�(���Y�ƅ�5��h"��<��u�u�%�e�o�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӖ��l^��G1�����u��
���L���YӖ��l_�'��&���������W��Y����G	�UךU���
�
�
�%�!�9�Mϗ�Y����)��tUךU���
�
�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�I����R��[
��U��������W�W���&ù��\��yN��1��������}�F�������V�=N��U���
�d�4�
�;�}�W���*����|!��d��Uʥ�e�d�u�u���3���>����v%��eN��@ʱ�"�!�u�|�]�}�W���&�ԓ�C9��SN�<����
���l�}�WϮ�I����	F��=��*����
����u�BϺ�����O��N�����d�
�%�#�3�g�>���-����t/��=N��U���
�a�o��w�	�(���0����p2��F�U���;�:�e�n�w�}����Hǹ��l��T��;ʆ�����]�}�W���&���/��d:��9�������w�l�W������]ǻN��*ڊ�`�4�
�9�w�}�9ύ�=����z%��N�����e�o�����;���:����g)��]����!�u�|�_�w�}�(ہ�&����_�!��U���
���n�w�}����H����f2��c*��:���
�����l��������l�N��A���4�
�9�u�w��W���&����p]ǻN��*ފ�u�u� �u���8���&����|4�_�����:�e�n�u�w�-�C�������WF��x;��&������_�w�}�(ہ�Y�ƃ�gF��s1��2������u�d�}�������9F���*ي�%�#�1�o��	�$���5����l�N��A��o������0���/����aF�N�����u�|�_�u�w��(ہ�	����\��b:��!�����n�u�w�-�C��Cө��5��h"��<������}�f�9� ���Y����F�G1��@���
�9�u�u��}�#���6����9F���*���u� �u����>���<����N��
�����e�n�u�u�'�i�A���&����	F��cN��1�����_�u�w��(���Y����`2��{!��6�����u�f�w�2����I��ƹF��hZ��*���#�1�o����3���>����F�G1��M��������4���:����U��S�����|�_�u�u���(������)��=��*����n�u�u�'�i�N��6����g"��x)��*�����}�d�3�*����P���F��1�����9�u�u� �w�	�(���0��ƹF��hZ��E��������4���:����U��S�����|�_�u�u���G���&����	F��cN��1�����_�u�w��(��Cө��5��h"��<������}�f�9� ���Y����F�G1��Dۊ�%�#�1�o��	�$���5����l�N��A��u�u� �u���8���&����|4�_�����:�e�n�u�w�-�C��&����_�!��U���
���n�w�}����H����|3��d:��9�������w�n�W������]ǻN��*ފ�f�4�
�9�w�}�"���-����t/��=N��U���
�a�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&�ғ�C9��SN�:��������W�W���&ǹ��\��b:��!�����
����_������\F��d��Uʥ�a�d�
�%�!�9�Mϑ�-ӵ��l*��~-�U���%�b�e�o��}�#���6����e#��x<��D���:�;�:�e�l�}�WϮ�N�֓�C9��SN�<����
���l�}�WϮ�N���/��d:��9�������w�l�W������]ǻN��*݊�
�%�#�1�m��W���&����p]ǻN��*݊�u�u�����0���/����aF�N�����u�|�_�u�w��(݁�	����\��yN��1�����_�u�w��(���Y����g"��x)��*�����}�`�3�*����P���F�� 1�����9�u�u����;���:���F�� 1�Oʜ�u��
����2���+������Y��E��u�u�%�b�c�<�(���Y�ƅ�5��h"��<��u�u�%�b�b�g�>���-����t/��a+��:���d�u�:�;�8�m�L���YӖ��lS��G1�����u��
���L���YӖ��lP�'��&���������W��Y����G	�UךU���
�
�
�%�!�9�Mϗ�Y����)��tUךU���
�
�u�u���3���>����v%��eN��@ʱ�"�!�u�|�]�}�W���&Ĺ��l��T��;ʆ�����]�}�W���&����z(��c*��:���
�����h��������l�N��B���4�
�9�u�w��$���5����l�N��B��o��u����>���<����N��
�����e�n�u�u�'�j�N���&����	F��=��*����n�u�u�'�j�F���Y����g"��x)��*�����}�`�3�*����P���F�� 1�*���#�1�o��w�	�(���0��ƹF��hY��D���u��
���(���-���S��X����n�u�u�%�`�l�(������/��d:��9����_�u�u���E��0�Ɵ�w9��p'��#����u�d�u�8�3���B�����h_�����9�u�u����;���:���F�� 1�U���������!���6���F��@ ��U���_�u�u�
��n��������z(��c*��:���n�u�u�%�`�l�W���7ӵ��l*��~-��0����}�`�1� �)�W���s���C9��Z�����1�o��u���8���B�����h_�Oʜ�u��
����2���+������Y��E��u�u�%�b�f���������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�
9��V�����u������4�ԜY�Ƽ�
9��N��U���
���
��	�%���Hӂ��]��G�U���%�l�d�4��1�W���7ӵ��l*��~-�U���%�l�g�o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�@�ԓ�C9��SN�<����
���l�}�WϮ�@���/��d:��9�������w�n�W������]ǻN��*ӊ�
�%�#�1�m��W���&����p]ǻN��*ӊ�u�u�����0���/����aF�N�����u�|�_�u�w��(ہ�	����\��yN��1�����_�u�w��(���Y����g"��x)��*�����}�d�3�*����P���F��1�����9�u�u����;���:���F��1�Oʜ�u��
����2���+������Y��E��u�u�%�l�a�<�(���Y�ƅ�5��h"��<��u�u�%�l�`�g�>���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��lQ��G1�����u��
���L���YӖ��l^�'��&���������W��Y����G	�UךU���
�
�
�%�!�9�Mϗ�Y����)��tUךU���
�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&ʹ��l��T��;ʆ�����]�}�W���&���/��d:��9�������w�n�W������]ǻN��*ӊ�e�4�
�9�w�}�9ύ�=����z%��N�����d�u�u����;���:����g)��]����!�u�|�_�w�}�(ց�H����E
��N��U���
���n�w�}����H����z(��c*��:���
�����l��������l�N��L��
�%�#�1�m��W���&����p]ǻN��*ӊ�f�o��u���8���&����|4�_�����:�e�n�u�w�-�N��&����_�'��&������_�w�}�(ց�M����}F��s1��2������u�d�}�������9F���*���4�
�9�u�w��$���5����l�N��L��u�u�����0���/����aF�N�����u�|�_�u�w��(�������WF��~ ��!�����u�n�2�9�}�������V��E�����u�3�8��n��2���Y���F�V�����0���
���6���7����|F��d:��;��u�u�4�!�>�(�ϝ�+����}#��c'��*����:�u�0�6�}�W�������G����U���w����b�;�Gö�
����V��hZ��=��������`����5����c3��q"��!��������/���I߮��l/��b:��4���-�b�e�e�;�i�C��1����}6��h-��6��`�e�e�e�{��(���,����p.��C��Ɲ�������E���L����.��h=��*���h�`�����#�������{*��d7��8���e������'��1����j(��qS�G����
��
��`�D���[���F��Y�����%�6�;�!�;�:���Cӵ��l*��~-��H��r�_�u�u�8�.��������]��[����o������M���I��ƹF��X �����4�
��&�f�;���Cӵ��l*��~-��0����}�u�:�9�2�G���D����V��UךU���:�&�4�!�6��#���I����9��Z1�Oʆ�������8���Lӂ��]��G��H���e�e�e�n�w�}��������R��c1��E���2�
�&�
�w�}�#���6����e#��x<��@ʱ�"�!�u�|�m�}�G��I����F�T�����u�%��
�'���������\��c*��:���
�����}�������	[�^�E���_�u�u�:�$�<�Ͽ�&����CV��C	�����a�o�����4���:����S��X����u�h�w�d�g�m�L���YӅ��@��CN��*���&�m�3�8�b�g�$���5����l0��c!��]���:�;�:�e�w�`�U��I���9F������!�4�
�:�$�����I����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�e�3�*����P���W�=N��U���&�4�!�4��2�����Г�\��c*��:���
�����h��������\�^�E��e�e�e�e�g�f�W�������R��V�����
�#�g�f�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�l�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Eʱ�"�!�u�|�m�}�G��Y����\��V �����:�&�
�#�e�i�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�F��B�����D��ʴ�
�:�&�
�!�o�F��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��H��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$��ځ�Y�Ɵ�w9��p'��#����u�a�1� �)�W���C���V��UךU���:�&�4�!�6�����&����lS�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��_�����u�:�&�4�#�<�(���
����9��T��!�����
����_�������V�S��D��e�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�d�w�]�}�W���
������T�����a�a�o����0���/����aF�
�����e�u�h�w�f�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Fʱ�"�!�u�|�m�}�G��[���F��Y�����%�6�;�!�;�i�O��*����|!��h8��!���}�u�:�;�8�m�W��[����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�f�3�*����P���W��L�U���6�;�!�;�w�-��������l%�=��*����
����u�W������F��L�E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Jӂ��]��G��H���e�e�n�u�w�>�����ƭ�l��D��ފ�u�u��
���(���-��� F��@ ��U���o�u�e�e�u�W�W�������]��G1�����9�a�f�o���;���:����g)��]�����:�e�u�h�u�m�F��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��I����F�T�����u�%�6�;�#�1�C��Cӵ��l*��~-��0����}�u�:�9�2�G���D����W�=N��U���&�4�!�4��2����ǹ��	F��s1��2������u�d�9� ���Y���F�^�N���u�6�;�!�9�}��������ER��T��!�����
����_�������V�S��D��w�_�u�u�8�.��������]��[��1��������4���Y����\��XN�U��w�d�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�g�m�L�ԜY�ƿ�T����6���&�u�u����>���<����N��S�����|�o�u�e�g�m�U�ԜY�ƭ�G��B�����0�6�1�;�w�}�������F��C�� ���3�8�0�6�3�3�W�������l ��T�����9�<�u�;�9��}���Y����R
��G1�����0�
��&�f�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�-�G�������TF��d:��9�������w�l�W������]ǻN�����9�%�e�e�'�8�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��w�_�u�u�>�3�Ϯ�I�֓�C9��S1��*���u�u��
���L���Yӕ��]��G1��E���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�m�F���&����	F��s1��2������u�f�}�������9F������%�e�d�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E���_�u�u�<�9�1����H����E
��^ �����u��
���f�W���
����_F��1�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�g�o��������`2��{!��6�����u�d�w�2����I��ƹF��^	��ʥ�e�g�%�0�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�W�ߊu�u�<�;�;�-�G�������W9��h��U����
���l�}�Wϭ�����C9��1��*���
�'�2�o���;���:���V�=N��U���;�9�%�e�d�4�(���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����f�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�����u�<�;�9�'�m�D���&����Z��^	��U���
���n�w�}�����Ƽ�9��V�����'�2�o����0���C���]ǻN�����9�%�e�a�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��E���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�g�i��������l��T��!�����n�u�w�.����Y����9��h��*���2�o�����4��Y���9F������%�e�`�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��@���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�e�b�<�(���&����Z�=��*����n�u�u�$�:����&ù��R��[
�����o������M���I��ƹF��^	��ʥ�e�c�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�e�c�6���������\��c*��:���n�u�u�&�0�<�W���&Ź��l��h���������g�W��B�����Y�����b�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9�� 1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�e�b�4��1�(���
���5��h"��<��u�u�&�2�6�}�(߁�&����_��E��Oʆ�����m�}�G��Y����Z��[N��E���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�e�m�4�
�;���������g"��x)��N���u�&�2�4�w��(ׁ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��L���
�<�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����
9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y�����l�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(�������A��N��1�����o�u�g�f�W���
����_F��1�*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�֓�9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y�����d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�m�F߁�	����l��PN�&������o�w�m�L���Yӕ��]��G1��Dۊ�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��lW��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�e�d�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G��&����_��E��Oʆ�����m�}�G��Y����Z��[N��E��
�;�&�2�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������lV��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�e�d�
�'�+����&����	F��s1��2���_�u�u�<�9�1����H����l��h���������g�W��B�����Y�����d�
�;�&�0�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������h_�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�e�d��-��������TF��d:��9����_�u�u�>�3�Ϯ�I����R��[
�����o������M���I��ƹF��^	��ʥ�e�d�
�;�$�:�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��h^��A���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�e�f���������@��N��1�����_�u�w�4����	�֓�9��h��*���2�o�����4��Y���9F������%�e�d�
�9�.���*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T����*���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�g�l�(�������]9��PN�&������_�w�}����Ӗ��lW��V�����'�2�o����0���C���]ǻN�����9�%�b�e�>�����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��B���%�0�u�u���8���&����|4�[�����:�e�u�h�u�m�G��I����V��UךU���<�;�9�%�`�m��������l��T��!�����n�u�w�.����Y����9��h��*���2�o�����4��Y���9F������%�b�d�<��4�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��D���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V�=N��U���;�9�%�b�f�<�(���&����Z�=��*����n�u�u�$�:����&Ĺ��R��[
�����o������M���I��ƹF��^	��ʥ�b�g�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F�� 1�����u�u��
���(���-���S��X����u�h�w�e�g�m�G��I����]ǻN�����9�%�b�g�6���������\��c*��:���n�u�u�&�0�<�W���&����l��h���������g�W��B�����Y�����f�<�
�<�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I���9F������%�b�f�4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�&����_��E��Oʆ�����m�}�G��Y����Z��[N��B���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�b�a�4�
�;���������g"��x)��N���u�&�2�4�w��(ہ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��@���
�<�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y�����`�4�
�9��3����Cӵ��l*��~-�U���&�2�4�u���(�������A��N��1�����o�u�g�f�W���
����_F�� 1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&Ĺ��C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��B���4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9�� 1��*���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&Ĺ��V�=��*����
����u�BϺ�����O�
N��E��e�e�e�e�g�m�L���Yӕ��]��G1��B���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(؁�&����\��c*��:���
�����h��������\�^�E��e�e�e�e�g�f�W���
����_F�� 1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����
9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(ց����5��h"��<������}�b�9� ���Y���F�^�E��e�e�e�e�l�}�Wϭ�����C9��1��*���
�;�&�2�m��3���>����F�D�����
�
�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����&Ĺ��l��D��Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�j�F߁����5��h"��<������}�b�9� ���Y���F�^�E��e�e�e�e�l�}�Wϭ�����C9��^�����1�<�
�<�w�}�#���6����9F������%�b�d�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����W��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�@��&����\��c*��:���
�����h��������\�^�E��e�e�e�e�g�f�W���
����_F�� 1�*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�b�d��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����H����V�=��*����
����u�BϺ�����O�
N��E��e�e�e�e�g�m�L���Yӕ��]��G1��D؊�%�#�1�<��4�W���-����t/��=N��U���;�9�%�b�f���������TF��d:��9����o�u�e�l�}�Wϭ�����C9��]�����2�o�����4���:����W��S�����|�_�u�u�>�3�Ϯ�N����C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��Y����Z��[N��B��
�%�#�1�>�����Y����)��tUךU���<�;�9�%�`�l�(�������A��N��1�����o�u�g�f�W���
����_F�� 1�*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ѓ�9��R	��U���
���
��	�%���Lӂ��]��G��H���e�e�e�e�g�m�G��B�����Y�����d�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�j�Fہ�	����l��PN�&������o�w�m�L���Yӕ��]��G1��Dߊ�;�&�2�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��lW��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I��ƹF��^	��ʥ�b�d�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�@��&����_��E��Oʆ�����m�}�G��Y����Z��[N��L���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�
9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ϯ�@�֓�C9��S1��*���u�u��
���L���Yӕ��]��G1��E���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�d�F���&����	F��s1��2������u�d�}�������9F������%�l�d�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ӊ�
�%�#�1�>�����Y����)��tUךU���<�;�9�%�n�l��������V�=��*����u�h�r�p�W�W���������h\�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�@�ԓ�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(݁�	����l��D��Oʆ�����]�}�W�������l_��h�����%�0�u�u���8���Y���A��N�����4�u�
�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ӊ�
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(ہ����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�l�c�<�(���&����Z�=��*����n�u�u�$�:����&ʹ��R��[
�����o������M���I��ƹF��^	��ʥ�l�`�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӗ��lS��G1�����
�<�u�u���8���B�����Y�����`�4�
�9��/���*����|!��T��R��_�u�u�<�9�1����O����@��N��1��������}�D�������V�=N��U���;�9�%�l�a�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����
�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�N�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*݊�;�&�2�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��lQ��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���&Ĺ��l��h�����o������}���Y����R
��hW��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u���(���
���5��h"��<������}�f�9� ���Y����F�D�����
�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L���4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
����������TF��d:��9����o�u�e�l�}�Wϭ�����C9��1��*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&ʹ��V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�d�N���&����Z��^	��U���
���n�w�}�����Ƽ�
9��V�����'�2�o����0���C���]ǻN�����9�%�l�d��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ӊ�e�%�0�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����R
��hW��E���
�9�
�;�$�:�Mύ�=����z%��N�����4�u�
�
�g�<�(���&����\��c*��:���u�h�r�r�]�}�W�������l_��1��*���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ד�A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(�������W9��h��U����
���l�}�Wϭ�����C9��_�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��o��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�l�d�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��L��
�%�#�1�>�����Y����)��tUךU���<�;�9�%�n�l�(�������A��N��1�����o�u�g�f�W���
����_F��1�*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ߓ� 9��R	��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�<�9�1����H����l��h�����o������}���Y����R
��hW��F���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�d�Fہ�����\��c*��:���
�����l��������l�N�����u�
�
�a�'�8�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��P ��U���
�a�4�
�;���������g"��x)��N���u�&�2�4�w��(�������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�
9��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����&ʹ��l��A�����<�u�u����>��Y����Z��[N��L��
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(ہ�����lW��E��C��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��1�����c�c�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�F ��E1�*؊�0�
�a�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��Q��*���`�'�2�c�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h�����d�
�
�0��j�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�a�l�%�:�A��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ފ� �3�'�d������I����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a�7�3�0��i�Fف�����F��d:��9�������w�n�W������]ǻN�����9�%�a�7�1�8�(���HŹ��T9�� N�&���������W��Y����G	�UךU���<�;�9�%�c�?����&�ғ�9��P1�E��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������S��1����f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����U��\��*���
�c�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��F���'�2�b�l�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lR��B����
�
�0�
�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�`�&�'�0�e�B��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������:�
�:�%�b�/���A����g"��x)��*�����}�u�8�3���B�����Y�����3�
�f�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hV�U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������`2��G^�����3�8�f�o���;���:���F��P ��U���&�2�7�1�b�m�MϜ�6����l�N�����u�%�'�2�'�4����	ù��F��d:��9����o�u�e�l�}�Wϭ�����V��T��D���2�g�f�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��@��T��*���%�e�&�2��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�:����&����CT�=��*����
����u�FϺ�����O��N�����4�u�0�
�c�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��*���$��
�%��)�G������5��h"��<��u�u�&�2�6�}��������lS��T��:����n�u�u�$�:����	����l��C�����<�d�o����0���C���]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�0�>�>��������9��T��!�����
����_�������V�=N��U���;�9�4�
�2�����&����P	��1����f�
�%�
�#�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��*���m�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��h��*��d�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	����T9��\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�ہ�����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�i����K����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�c�1��@܁�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�0��m�F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����
� �m�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��M���2�g�b�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��R	��E��o������!���6�����Y��E��u�u�&�2�6�}�����Փ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����V��T��!�����
����_�������V�=N��U���;�9�3�
�#���������lV��_�� ��`�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��_��X�����d�
�
�=��8�(��M����g"��x)��*�����}�d�3�*����P���F��P ��U���-� �,� �����Oƹ��\��c*��:���
�����h��������l�N�����u��-� �.�(�(�������_�=��*����
����u�BϺ�����O��N�����4�u�0�
�:�l�(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����K����	F��s1��2������u�g�9� ���Y����F�D�����%�'�2�%�$�:��������l��h\�A���e�<�d�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��*��`�o�����4���:����V��X����n�u�u�&�0�<�W�������C��h��*���d�
�0�
�f�h�������5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�`�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���
�%�!�
�2����&����W��h��*���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}��������A��_�U����
�����#���Q�ƨ�D��^����u�<�;�9�6�����	����@��C��C���2�g�a�
�'�����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
� �d�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����b�'�2�g�b�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������E�����2�&�9�!�'�j����K����C��^�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������S��N��1��������}�GϺ�����O��N�����4�u�%�'�0�-����
����^��h��*��l�%�e�<�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��L���
�d�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���
�d�`�o���;���:����g)��^�����:�e�n�u�w�.����Y����V��G��*���
�8�d�
�2��F���	�֓�GW�=��*����
����u�W������]ǻN�����9�3�
�!��/�;���&�ғ�l��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"����
�
�=�
�2��F��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��"��� �,� �
�`�l����K�ѓ�F��d:��9�������w�l�W������]ǻN�����9�<�
������&¹��T9��\��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u��1�(���&����lS��h_�� ��l�
�g�o���;���:����g)��Z�����:�e�n�u�w�.����Y����Z9��E1�����
�
�
�0��l�@��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Q=�����!�'�
�
�"�l�Nց�H����g"��x)��*�����}�d�3�*����P���F��P ��U���&�2�6�0��	����
����U��N�&������_�w�}����Ӈ��@��U
��M��o�����W�W������� ��Y��*���8�a�
�
�"�l�G܁�H����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �3�'�f��(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
�"�;���&¹��T9��\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u����������9��h_�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��1�����g�e�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��A���3�
�f�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�a�m�'�0�o�F���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���3�0�
�a�f����Nù��\��c*��:���
�����l��������l�N�����u�
�
� �1�/�Fہ�J����lT�� N�&���������W��Y����G	�UךU���<�;�9�%�c�?����&�ғ�9��h_�@���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����V��1�*���
�g�g�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��Q��Dފ�b�3�
�a�`�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�a�g��8�(��N����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �3�'�f��C���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����M����A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�F ��E1�*���'�2�g�f�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��U�����`�d�3�
�b�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��A���3�0�
�`�f�/���M����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a�7�3�0��h�C���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����L�ғ�V��Z�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�i��������l^��B1�M݊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����U��[��*���
�g�g�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��Q��Dߊ�f�3�
�c�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�`�d��8�(��N����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �3�'�f��F���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����L����U��W�����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����lW��Z�� ��a�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��Q��Dߊ�d�3�
�b�g�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^"�����'��:�
��5�(���A�ԓ�F��d:��9�������w�i��������l�N�����u�%�&�2�4�8�(���
�ޓ�@��T��!�����n�u�w�.����Y����Z��S
��D���u����l�}�Wϭ�����T��Q��Gӊ�e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����U��G^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:����H����	F��s1��2������u�d�9� ���Y����F�D�����'�6�;�
�"�d�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����9�3�
�l��n�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��R��ۊ� �l�l�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����\��X ��*���l�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӊ��P	��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/����J����
R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;� �8�C���&����CU�=��*����
����u�BϺ�����O��N�����4�u�0��;����J����	F��s1��2������u�f�}�������9F������;�"�0�b�1��Aց�J����g"��x)��*�����}�`�3�*����P���F��P ��U����9�
� �n�h����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����l�3�
�m��n�Mύ�=����z%��r-��'���`�1�"�!�w�t�}���Y����R
��R�����3�
�m�
�d�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������d��D���
�l�
�f�m��3���>����v%��eN��@ʱ�"�!�u�|�]�}�W�������V��[_�����e�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��G[�� ��d�
�f�o���;���:����g)��]����!�u�|�_�w�}����ӕ��l�� 1��*��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��h��D���
�f�o����0���/����aF�N�����u�|�_�u�w�4��������_P��B1�D���u�u��
���(���-���S��X����n�u�u�&�0�<�W���*����l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l*��G1��D��e�!�3�
�g�l����Y����)��t1��6���u�f�1�"�#�}�^�ԜY�ƿ�T�������m�3�
�d�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����3�
�d�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��@=��Dߊ� �d�f�
�d�g�$���5����l0��c!��]���1�"�!�u�~�W�W�������	��T��L���
�d�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A9��Y
�����d�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӈ��`��1��*��f�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����V
��h��D���
�f�o����0���/����aF�N�����u�|�_�u�w�4��������]��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����9��h_�D���u�u��
���(���-���S��X����n�u�u�&�0�<�W���*����l ��_�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������U��W�����u��
����2���+������Y��E��u�u�&�2�6�}�����ԓ�F9��Y��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���K����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���M����T��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*���&����W��G]��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u�2���������U��N�&���������W��Y����G	�UךU���<�;�9�&�;�)�������� _��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������S��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������T��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������_��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������P��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������U��N�&���������W��Y����G	�UךU���<�;�9�;� �8�E߁����� 9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��1�@���&����l��N��1��������}�F�������V�=N��U���;�9�%�a�5�;����M�Փ�F9��Z��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������R��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�F ��E1�*݊� �d�f�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h�����d�
�e�3��n�N���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����7�3�0�
�c�l�(���H����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
�"�;���&�ԓ�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������R�� 1��*��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��A��
� �d�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hZ�� ���'�d�
�l�1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a�7�3�0��i�E߁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�
��(����Hǹ��l ��Z�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��h\�����a�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��Q��*���g�
� �d�e��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�'�d�
�b�;�(��J����	F��s1��2������u�d�}�������9F������%�a�7�3�2��C��&����R��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u����������^��B1�@ފ�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����U��Z��L���
�a�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��U�����a�f�
� �f�k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ފ� �3�'�d��l����M�ӓ� F��d:��9�������w�n�W������]ǻN�����9�%�a�7�1�8�(���J����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�F ��E1�*���3�
�`�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�a�f�
�"�l�F߁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �3�'�f��@���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����M����U��\�����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����lW��W�� ��f�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��Q��Dފ�e�3�
�`�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�`�f�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a�7�3�0��h�A���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����L�ѓ�F9��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�C�������S��1��*���a�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��@��
� �d�e��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hZ�� ���'�d�
�g�1��A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�a�7�3�0��h�F؁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�
��(����Hƹ��l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��h_�����c�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��Q��*���g�
� �d�c��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�'�d�
�e�;�(��N����	F��s1��2������u�d�}�������9F������%�a�7�3�2��B��&����P��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u����������R��B1�Bۊ�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�M����U��[��@���
�c�m�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��U�����`�g�
� �f�e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ފ� �3�'�d��e����O�ߓ� F��d:��9�������w�n�W������]ǻN�����9�%�a�7�1�8�(���Kʹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ғ�F ��E1�*���3�
�b�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�`�f�
�"�l�E؁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �3�'�f��D���&����l��N��1��������}�D�������V�=N��U���;�9�%�a�5�;����L����U�� Z�����u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����lW��X�� ��`�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��Q��Dߊ�b�3�
�b�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�`�f��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����
�
� �3�%�l�(�������P��N�&���������W��Y����G	�UךU���<�;�9�%�c�?����&�ӓ�9��h_�F���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&���� U��RN�&������_�w�}����Ӈ��}5��D��U���
���
��	�%���Y����G	�UךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����P��T��:����n�u�u�$�:����	����l��hW�U������n�w�}�����ƭ�l��h��*��o�����W�W���������D�����d�d�o����9�ԜY�ƿ�T�������7�1�d�e�m��8���7���F��P ��U���&�2�7�1�f�d�MϜ�6����l�N�����u�%�&�2�5�9�F��CӤ��#��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w�-��������P�,��9���n�u�u�&�0�<�W���
����W��N�7�����_�u�w�4��������T9��S1�U������n�w�}�����ƭ�l��h��*��o�����W�W���������D�����b�u�u����L���Yӕ��]��V�����1�
�c�o���2���s���@��V�����2�7�1�l�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��m�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�<�(���&����W��N��:����_�u�u�>�3�Ͽ�&����Q��^�Oʗ����_�w�}����Ӈ��@��U
��F��o�����W�W���������D�����f�`�o����9�ԜY�ƿ�T�������7�1�f�a�m��8���7���F��P ��U���&�2�7�1�d�n�MϜ�6����l�N�����u�%�&�2�5�9�D��CӤ��#��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-�������� S�,��9���n�u�u�&�0�<�W���
����W��Z��U�����n�u�w�.����Y����Z��S
��@���u����l�}�Wϭ�����R��^	�����c�u�u����L���Yӕ��]��V�����1�
�b�u�w��;���B�����Y�����<�
�1�
�o�}�W���5����9F������4�
�<�
�3��O���Y����v'��=N��U���;�9�4�
�>�����@����q)��r/�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��S1�E������]�}�W�������C9��P1����l�o�����}���Y����R
��G1�����1�a�m�o���2���s���@��V�����2�7�1�a�`�g�5���<����F�D�����%�&�2�7�3�i�A��;����r(��N�����4�u�%�&�0�?���I����|)��v �U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������lU��T��:����n�u�u�$�:����	����l��h]�U������n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���
�d�u�u���6��Y����Z��[N��*���
�1�
�g�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��n�W���6����}]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUװU���6�8�:�0�#�0�6���8ƣ��9��B��G���f�;�
�g�f�0����	ӯ��F�P�����}�u�u�u�w��W���7����a]ǻN��U��� �
���w�}�9���<��ƹF�N��������o��	�0���s���F�S��*����u�u����L���Y�����C1��1���o�����t�}���Y����NǻN��U���<�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������	F��=��*����
����u�FϺ�����O��N��U���1� �u�u��}�#���6����e#��x<��F���:�;�:�e�w�f�W�������\��Y��N�ߠu�u�6�8�8�8�ϳ�8�߈�#��1�����
�g�
�g�e��}���Y����A��d��U���u��u�u���2��Y���F��b#��!���u�u����f�W���Y����Z��`'��=������]�}�W���Y����l1��c&��U�����u�n�w�}����Y���F�N�����u��
���L���Y�����R��U��������W�W���Y�ƨ�]V�'��&���������W��Y����G	�UךU���u�u�0�o��}�#���6����9F�N��U���!�o�����;���:����g)��]����!�u�|�|�]�}�W���Y����\��CUװ��2�;�u�u�1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�
�g�g����������vW��@���e�3� �
�e�.�Dݰ�&�ԓ�l��h
�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��|�u�u�%�%�}����s���F�S��U��2�%�3�
�e��G�ԜY���F��Y_��Kʧ�2�m�c�_�w�}�W������F��G1��*��
�g�n�_�w�}�(߁�����lU��h]��G���u�u�:�%�9�3�W���8ʢ��v ��h�����f�&�f�
�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�:�!� ��?��Y���F�G��U���u�_�u�u�w�}����GӇ��P
��=N��U���u�0�0�u�i�<�(���U���F�
��E��u�'�
� �o�n���Y���F��RN��U���
� �m�f�4�q�W���Y����\��
P����� �m�f�%�~�W�}�ԶY���F��RN�����!�&�4�0��-�4���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�_�u�u�w�}�W���Y���F��h-�����i�u�%���.�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�4�
�0��-����	�֓�GV��D��ʥ�:�0�&�u�z�}�WϿ�&����C��R ��ڊ�!�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}��������G��G����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}��������T9��S1�G���!�0�u�u�w�}�W���Y���F�N��U���'�2�%�<�2��߁������T�����2�6�e�_�w�}�W���Y���F�N�����}�%�&�2�5�9�A��Y����l�N��U���u�u�u�u�w�}�WϿ�&����C��R ��ڊ�!�u�h�4��2��������]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u�'�/��������C��^����2�u�'�6�$�s�Z�ԜY�ƭ�l��h�����%�e�<�d�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W�������T9��^��*���
�!�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���!�:�1�
�2��G��DӇ��P	��C1��D��u�;�u�4��2��������F�V�����&�$��
�'���������O�C��U���u�u�u�u�w�}�W���YӇ��A��G�����%�
�!�u�j�<�(���
����T��UךU���u�u�u�u�w�}����Y���R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1��\ʴ�1�;�!�4��4�(���&����F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��E���2�
�&�
�~�<�ϰ��Ω�Z��Y
�����g�f�u�u�'�>�����ד�O�N�����u�u�u�u�w�}�W���Y����C9��P1�����
�%�
�!�w�`��������_	��T1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lV��G1�����0�u�&�<�9�-����
���9F���*ڊ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�e�e�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��l�W������F�N��U���u�u�u�u�w�-�G�������W9��R	��Hʥ�e�e�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ڊ�
�'�2�4�$�:�W�������K��N�����e�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�
�
��-����Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�~�}����s���F�N��U���u�u�%�e�g�-����DӖ��lV��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&�֓�C9��S1�����&�<�;�%�8�8����T�����h_�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�9��h��*���2�i�u�%�4�3��������l�N��U���u�0�&�_�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&�����Yd��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�$�:����&����G^��D��\���=�;�_�u�w�}�W���Y���F�N�����d�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�f�l�W������F�N��U���u�u�u�u�w�-�G��&����_��E��I���
�
�e�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�e�%�0�w�.����	����@�CךU���
�
�e�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e�d�
�'�+����Y����l�N��U���u�u�u�u�w�-�G��&����Z�G1��D��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��_�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�d�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^��D���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:��Ҋ�&�
�|�u�?�3�}���Y���F�N��U���u�u�%�e�f���������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����H���G��d��U���u�u�u�u�w�}�W���YӖ��lW��V�����'�2�i�u���F���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��l����Y����T��E�����x�_�u�u���F�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��E��
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m�Fށ�	����O�C��U���u�u�u�u�w�}�W���YӖ��lW��G��U��%�e�d�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����d�
�%�#�3�-����
������T��[���_�u�u�
��o��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�g�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���u�u�u�u�w�}����H����l��h����u�%�6�;�#�1����I���F�N��U���u�u�u�0�$�;�_���
����W��W�����u�u�u�u�w�}�W���Y���F���*���4�
�9�
�%�:�K���&ù��l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&�ԓ�A��V�����'�6�&�{�z�W�W���&ù��l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�e�d��/���Y����\��h��C��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�֓�9��h��\���!�0�u�u�w�}�W���Y���F���*���%�0�u�h�'�m�F��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�e�f���������TF��D��U���6�&�{�x�]�}�W���&�Փ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���D���&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��<�(���
����T��N�����<�
�&�$���ׁ�
����F��R ��U���u�u�u�u�w�}�W���Y����lV��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����`�|�!�0�w�}�W���Y���F�N��U���u�
�
�f�6��������F��1�*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��]�����4�&�2�u�%�>���T���F��1�*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G��&����Z�V�����
�#�c�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h^��F���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�f�'�8�W��	�֓� ]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����Hǹ��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��Z�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��l��A�����u�h�4�
�8�.�(�������9F�N��U���u�9�0�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ڊ�a�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�a�t����Y���F�N��U���u�u�u�u�w��(�������W9��R	��Hʥ�e�d�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����d�
�'�2�6�.��������@H�d��Uʥ�e�d�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lW��G��U��4�
�:�&��+�A��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�a�4��1�^�������9F�N��U���u�u�u�u�w��(���	����[��h^��A�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��1��*���
�'�2�4�$�:�W�������K��N�����d�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��M���8�`�|�!�2�}�W���Y���F�N��U���u�u�
�
�b�<�(���&����Z�V�����
�:�<�
�l�}�W���Y���F�N��U���<�u�4�
�>�����N����[��=N��U���u�u�u�u�w�}�W���Y����S��G1�����0�u�h�%�g�l�(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�e�f���������]F��X�����x�u�u�%�g�l�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���B���&����O��_�����u�u�u�u�w�}�W���Y����S��E��I���
�
�`�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ڊ�
�%�#�1�'�8�W�������A	��D�X�ߊu�u�
�
��-����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����d�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N��U���u�u�u�u�'�m�F���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lV��h�����%�0�u�h�'�m�F���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�g�l����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��D���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�I�ד�A��S��*ڊ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����9�
�'�2�6�.��������@H�d��Uʥ�e�g�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��M���8�`�|�!�2�}�W���Y���F�N��U���u�u�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���PӒ��]FǻN��U���u�u�u�u�w�}�W���&ù��R��[
�����i�u�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�e�g�%�2�}����Ӗ��P��N����u�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lV��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�e�g�4��1�^�������9F�N��U���u�u�u�u�w��(݁����F��1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lU��G1�����0�u�&�<�9�-����
���9F���*ي�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�e�f�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��e�W������F�N��U���u�u�u�u�w�-�G�������W9��R	��Hʥ�e�f�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ڊ�
�'�2�4�$�:�W�������K��N�����f�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��C��R�����:�&�
�#�a�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ڊ�
�%�#�1�~�}����s���F�N��U���u�u�%�e�d�-����DӖ��lU��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&ǹ��l��h��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�I�ғ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�W���Y���F���*ފ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�b�|�#�8�W���Y���F�N��U���u�u�u�
����������TF���*ފ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����u�&�<�;�'�2����Y��ƹF��h^��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�-�G���	����[��G1�����9�d�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�|�!�2�}�W���Y���F�N��U���
�
�
�'�0�a�W���&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�B���&����C�������%�:�0�&�w�p�W���	�֓�l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(ځ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�}�W���Y���C9��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����c�u�=�;�]�}�W���Y���F�N��U���%�e�`�4��1�(������C9��1��*���n�u�u�u�w�}�W���Y����������u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lS��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��lS��G1�����u�=�;�_�w�}�W���Y���F�N��E���%�0�u�h�'�m�B�ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��-����	����R��P �����&�{�x�_�w�}�(߁�&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�e�a�<�(���&����Z�V�����
�:�<�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�u�u�w�}�W���	�֓�l��A�����u�h�4�
�8�.�(�������9F�N��U���u�u�u�u�w�1��������T9��S1�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ڊ�
�%�#�1�'�8�W��	�֓�l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&Ź��V��D��ʥ�:�0�&�u�z�}�WϮ�I�Г�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e�c�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&Ź��l��G�����u�u�u�u�w�}�W���Y�����hX�����i�u�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�e�b�4�
�;���������]F��X�����x�u�u�%�g�j��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�m�3�:�h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lW��N�����u�u�u�u�w�}�W���Y���F��h^��*���#�1�%�0�w�`����N����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(؁�����@��YN�����&�u�x�u�w�-�G���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����b�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(؁�	����O�C��U���u�u�u�u�w�}�W���YӖ��lQ��E��I���
�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��E���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�e�m�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���m�3�8�`�~�)����Y���F�N��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lV��h�����%�0�u�h�'�m�O���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�g�e����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��M���0�u�h�4��2�����Г�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�I�ޓ�A��S��*ڊ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����9�
�'�2�6�.��������@H�d��Uʥ�e�l�4�
�;���������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h^��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��M���8�`�|�!�2�}�W���Y���F�N��U���u�u�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���K�Ƹ�V�N��U���u�u�u�u�w�}�W���	�֓�l��A�����u�h�%�e�n�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
�%�:�����Ƽ�\��D@��X���u�%�e�l�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�
�'�+����Y����l�N��U���u�u�u�u�w�-�G���	����[��h^��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��V�����'�2�4�&�0�}����
���l�N��B���4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��h�����%�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y�����T�����2�6�d�h�6�����
����g9��1�����|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�o�@������F�N��U���u�u�u�u�w�}����I����E
��G��U��%�b�e�4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�'�2�6�.��������@H�d��Uʥ�b�e�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����9��R	��Hʴ�
�:�&�
�!�k�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�W������F�N��U���u�u�u�%�`�m����Y����lQ��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��l��A�����u�&�<�;�'�2����Y��ƹF��hY��E���
�9�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��lW��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�b�d�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y���F�R�����%�&�2�7�3�n�@������F�N��U���u�u�u�u�w�}����Hù��l��h����u�
�
�e�6����Y���F�N��U���u�u�;�u�1�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�e�%�2�}����Ӗ��P��N����u�
�
�e�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��^�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�b�d��-����P�Ƹ�V�N��U���u�u�u�u�w�}����Hù��V�
N��B��n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�*���#�1�%�0�w�.����	����@�CךU���
�
�d�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N��U���u�u�u�%�`�l�(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����lQ��1��*���
�'�2�i�w��(�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���F����ƭ�@�������{�x�_�u�w��(���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����d�
�'�2�k�}��������EW��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@��&����_�N�����u�u�u�u�w�}�W���Y����lQ��1�����h�%�b�d�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b�d�
�%�!�9����Y����T��E�����x�_�u�u���E���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�g�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�u�u�u�w�}�WϮ�N����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h]�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�g�4�
�9��/���Y����T��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&Ĺ��l��PN�����u�'�6�&�y�p�}���Y����T��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b�f�����E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��lW��V�����|�!�0�u�w�}�W���Y���F�N��*݊�g�%�0�u�j�-�@��B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`�l�(�������A��V�����'�6�&�{�z�W�W���&Ĺ��l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�}�W���Y�����h_�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
�d�<�(���&����Z�G1��Dي�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F�� 1�*���2�4�&�2�w�/����W���F�G1��Dي�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����H����V�
N��*���&�
�#�c�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�
�9�|�~�)����Y���F�N��U���u�u�
�
�d�-����DӖ��lW��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�N����R��[
�����4�&�2�u�%�>���T���F�� 1�*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����R��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��Q��@���!�0�u�u�w�}�W���Y���F�N��U���
�a�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��i�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�M����E
��G��U��%�b�d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b�d�
�'�0�<����Y����V��C�U���%�b�d�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�a�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(؁�M����TF���*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h_�����9�
�'�2�6�.��������@H�d��Uʥ�b�d�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��Dߊ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
��h��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��h�����%�0�u�h�'�j�Fځ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`�l�(���Ӈ��Z��G�����u�x�u�u�'�j�Fځ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�`�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�9��h����u�
�
�`�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�%�#�3�-����
������T��[���_�u�u�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�b�d�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��U���u�u�u�u�w�-�@�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����T�����ߊu�u�u�u�w�}�W���Y���F�� 1�����9�
�'�2�k�}�(؁�&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�j�F����ƭ�@�������{�x�_�u�w��(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*݊�
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�j�F���&����O��_�����u�u�u�u�w�}�W���Y����9��R	��Hʥ�b�d�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*؊�%�#�1�%�2�}����Ӗ��P��N����u�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��B���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N��U���u�u�u�%�`�o��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b�e�-����
������T��[���_�u�u�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hY��*���2�i�u�%�4�3����HŹ��9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�b�e�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����V�
N��B��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h]�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F�N��U���u�%�b�f�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��R��[
�����i�u�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�b�f�%�2�}����Ӗ��P��N����u�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lQ��h����u�%�6�;�#�1�Fف�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�b�f�4��1�^�������9F�N��U���u�u�u�u�w��(܁����F�� 1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lR��G1�����0�u�&�<�9�-����
���9F���*ފ�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�b�a�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&����_��E��I���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����a�%�0�u�$�4�Ϯ�����F�=N��U���
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ѓ�l��PN�U���6�;�!�9�f��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����a�4�
�9�~�t����Y���F�N��U���u�u�u�
������E�Ƽ�9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�N�ӓ�C9��S1�����&�<�;�%�8�8����T�����h[�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&Ĺ��R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����l ��h[��U���;�_�u�u�w�}�W���Y���F�N��B���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�c�~�)����Y���F�N��U���u�u�u�u���(�������A��S��*݊�
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��@���0�u�&�<�9�-����
���9F���*ߊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����L����TF������!�9�d�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��@���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�
�%�:�K���&Ĺ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�@�������W9��R	�����;�%�:�0�$�}�Z���YӖ��lP��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(؁�&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���A����lS����ߊu�u�u�u�w�}�W���Y���F�� 1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�b�|�!�2�}�W���Y���F�N��U���u�u�
�
��-����	����[��hY��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��1�����&�<�;�%�8�8����T�����hX�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�j�A��������T�����d�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�'�2�k�}�(؁�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�`�j��������V��D��ʥ�:�0�&�u�z�}�WϮ�N�ѓ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�O��������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����lQ��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����9��R	�����;�%�:�0�$�}�Z���YӖ��lQ��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�b�`�-����DӇ��P	��C1��D܊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����9��h��\���!�0�u�u�w�}�W���Y���F���*݊�'�2�i�u���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�b�m�6���������@��YN�����&�u�x�u�w�-�@�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�o�;���PӒ��]FǻN��U���u�u�u�u�w�}�W���&Ĺ��R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��h\�\ʡ�0�u�u�u�w�}�W���Y���F�N��*݊�
�%�#�1�'�8�W��	�ѓ�l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&˹��V��D��ʥ�:�0�&�u�z�}�WϮ�N�ޓ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�b�m�%�2�}�JϿ�&����G9��X��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&˹��l��G�����u�u�u�u�w�}�W���Y�����hV�����i�u�
�
�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�b�l�4�
�;���������]F��X�����x�u�u�%�`�d��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�m�3�:�h�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(؁�&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lT��N�����u�u�u�u�w�}�W���Y���F��hY��*���#�1�%�0�w�`����@����E
��=N��U���u�u�u�u�w�}�W���Y����F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w��(ց�����@��YN�����&�u�x�u�w�-�@���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����l�%�0�u�j�<�(���
����P��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(ց�	����O�C��U���u�u�u�u�w�}�W���YӖ��l_��E��I���
�
�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��L���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�l�e�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ӊ�
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^��]���6�;�!�9�0�>�F������T9��R��!���m�3�8�`�~�)����Y���F�N��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����l_��h�����%�0�u�h�'�d�G���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�n�m����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��E���0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�@�֓�A��S��*ӊ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�*���#�1�%�0�w�.����	����@�CךU���
�
�e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N��U���u�u�u�%�n�l�(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.��������F��R ��U���u�u�u�u�w�}�W���Y����l_��1��*���
�'�2�i�w��(�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���G����ƭ�@�������{�x�_�u�w��(���	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����d�
�'�2�k�}��������EU��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�N��&����_�N�����u�u�u�u�w�}�W���Y����l_��1�����h�%�l�d�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�l�d�
�%�!�9����Y����T��E�����x�_�u�u���F���&����C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�d�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�u�u�u�w�}�WϮ�@����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hZ�\ʡ�0�u�u�u�w�}�W���Y���F�N��*ӊ�d�4�
�9��/���Y����W��G1���ߊu�u�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&ʹ��l��PN�����u�'�6�&�y�p�}���Y����W��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l�f�����E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��lW��V�����|�!�0�u�w�}�W���Y���F�N��*ӊ�d�%�0�u�j�-�N��B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�n�l�(�������A��V�����'�6�&�{�z�W�W���&ʹ��l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�}�W���Y�����h_�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�c�|�!�2�}�W���Y���F�N��U���u�u�
�
�e�<�(���&����Z�G1��D؊�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�*���2�4�&�2�w�/����W���F�G1��D؊�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����H����V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�
�9�|�~�)����Y���F�N��U���u�u�
�
�e�-����DӖ��lW��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�@����R��[
�����4�&�2�u�%�>���T���F��1�*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����U��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��Q��@���!�0�u�u�w�}�W���Y���F�N��U���
�f�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��j�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ց�J����E
��G��U��%�l�d�
�'�+��ԜY���F�N��U���u�0�1�<�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʥ�l�d�
�'�0�<����Y����V��C�U���%�l�d�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����l_��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�f�6�����PӒ��]FǻN��U���u�u�u�u�w�}�(ց�J����TF���*��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h_�����9�
�'�2�6�.��������@H�d��Uʥ�l�d�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��Dފ�%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�#�8�W���Y���F�N��U���u�u�u�
��i��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�
9��h�����%�0�u�h�'�d�Fہ�	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�n�l�(���Ӈ��Z��G�����u�x�u�u�'�d�Fہ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ӊ�a�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������WO����ߊu�u�u�u�w�}�W���Y�Ƽ�
9��h����u�
�
�a�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�`�4�
�;���������]F��X�����x�u�u�%�n�l�(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�l�d�
�'�+���������T�����2�6�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�W�W���Y���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�m�1�0�B�������9F�N��U���u�u�u�u�w�}�W���&�ӓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��W�U���;�_�u�u�w�}�W���Y���F�N��L��
�%�#�1�'�8�W��	�ߓ�9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�@����C�������%�:�0�&�w�p�W���	�ߓ�9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�b�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����S��G1�����u�=�;�_�w�}�W���Y���F�N��L��
�'�2�i�w��(��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������TF��D��U���6�&�{�x�]�}�W���&¹��l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�n�l��������V�
N��*���&�
�:�<��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��lW��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��F��u�=�;�_�w�}�W���Y���F�N��Uʥ�l�d�4�
�;�����E�Ƽ�
9��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�l��PN�����u�'�6�&�y�p�}���Y����9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ�l��A��\���=�;�_�u�w�}�W���Y���F�G1��D���0�u�h�%�n�l�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�
�'�+�����ƭ�@�������{�x�_�u�w��(݁�	����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�l�g�6��������F��h�����:�<�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�u�u�u�w�}�WϮ�@�ԓ�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��Y�U���;�_�u�u�w�}�W���Y���F�N��L���4�
�9�
�%�:�K���&ʹ��R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����K����TF��D��U���6�&�{�x�]�}�W���&����V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`����K����E
��G�����_�u�u�u�w�}�W���Y���C9��1�����h�%�l�g�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�%�#�3�-����
������T��[���_�u�u�
����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�l�f�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��U���u�u�u�u�w�-�N�������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&���� ^�����ߊu�u�u�u�w�}�W���Y���F��1�����9�
�'�2�k�}�(ց�&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�d�D����ƭ�@�������{�x�_�u�w��(܁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ӊ�
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�d�D���&����O��_�����u�u�u�u�w�}�W���Y���� 9��R	��Hʥ�l�f�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*ފ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��L���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N��U���u�u�u�%�n�i��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&������YNךU���u�u�u�u�w�}�W���Y�Ƽ�
9��V�����'�2�i�u���(�������F�N��U���u�u�u�u�2�9���Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�l�c�-����
������T��[���_�u�u�
����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��hW��*���2�i�u�%�4�3����J����9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�l�c�<�(���P����[��=N��U���u�u�u�u�w�}�W���&ǹ��V�
N��L��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����h[�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�
�%�#�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F�N��U���u�%�l�`�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�W���&ʹ��R��[
�����i�u�
�
��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�l�`�%�2�}����Ӗ��P��N����u�
�
�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����l_��h����u�%�6�;�#�1�D݁�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�l�`�4��1�^�������9F�N��U���u�u�u�u�w��(ځ����F��1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��lP��G1�����0�u�&�<�9�-����
���9F���*܊�%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�
9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��*���u�=�;�_�w�}�W���Y���F�N��Uʥ�l�c�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W���Y���F��[��U´�
�<�
�1��l�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ց�&����_��E��I���
�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����c�%�0�u�$�4�Ϯ�����F�=N��U���
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ߓ�l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����c�4�
�9�~�t����Y���F�N��U���u�u�u�
������E�Ƽ�
9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�@�ѓ�C9��S1�����&�<�;�%�8�8����T�����hY�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ʹ��R��[
�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����l ��h[��U���;�_�u�u�w�}�W���Y���F�N��L���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�g�~�)����Y���F�N��U���u�u�u�u���(�������A��S��*ӊ�
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��B���0�u�&�<�9�-����
���9F���*݊�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����N����TF������!�9�f�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��B���
�9�|�|�#�8�W���Y���F�N��U���u�
�
�
�%�:�K���&ʹ��9F�N��U���u�u�u�;�w�;�W���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�_�u�u�z�-�N�������W9��R	�����;�%�:�0�$�}�Z���YӖ��l^��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ց�&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���A����lS����ߊu�u�u�u�w�}�W���Y���F��1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�w�}�W�������N��h��*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
��-����	����[��hW��*���#�1�_�u�w�}�W���Y���F�R ����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��1�����&�<�;�%�8�8����T�����hV�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�d�O��������T�����f�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�
�'�2�k�}�(ց�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�n�d��������V��D��ʥ�:�0�&�u�z�}�WϮ�@�ߓ�C9��S1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�O��������YNךU���u�u�u�u�w�}�W���Y�Ƽ�
9��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�
�%�!�9����Y����l_��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����
9��R	�����;�%�:�0�$�}�Z���YӖ��l_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�l�n�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����
9��h��\���!�0�u�u�w�}�W���Y���F���*ӊ�'�2�i�u���L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�<�
�<��/�;���&ƹ��T9��N�����u�'�6�&�y�p�}���Y����Z9��E1�����
�0�
�d��.����	����	F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�u�u�w�}�;���&����	��h[�����d�u�h�<��4�1���5����9��1����m�n�u�u�w�}�W���Y����_��F��*���
�1�
�b�~�)����Y���F�N��U���u�u��9��2�(���	�ӓ�V��V��Hʴ�
�:�&�
�!��L���Y���F�N��U���u�3�_�u�w�}�W���Y����Z ��=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����@��h��*���|�!�0�_�w�}�W���Y���F��h��*���!�
�-�!�8�9�(���&����l��h��U��0�<�6�;�f�/���J��ƹF�N��U���u�u�%�'�0�-����
����^��h��*��a�%�e�<�f�a�W���&���� 9��P1�D��u�u�u�u�w�}�W�������T9��D�����!�%�a�'�0�o�Eځ�	ù��F���*���d�
�0�
�f�h�}���Y���F�N�����0�
�%�!��8�(���Hƹ��T9��[��ڊ�!�u�h�&�;�)��������U��=N��U���u�u�u�u�w�-����	����l��h��D܊�0�
�d�a�'�m���E�ƿ�_9��G_�����g�a�n�u�w�}�W���Y�����E�����2�&�9�!�'�j����K����C��^�I���0�
�8�d��8�(��K���F�N��U���u�4�
�0��-��������CW��E��G���
�%�
�!�w�`��������l��h\�L�ߊu�u�u�u�w�}�W���	����l��C	�����8�d�
�0��l�B���I����Z�D�����l�'�2�g�a�f�W���Y���F�N�����:�1�
�0��m�@��Y����P	��1��*��
�g�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���	�֓�G��Q��D���;�u�4�
�8�.�(���&���V��T��D���
�a�
�g�~�}����Y���F�N��U����9�
�:��2���&ù��Z9��P1�E���h�3�
�!��/�;���&�ғ�l��h��D���
�f�_�u�w�}�W���Y���U5��C1�����:�
�a�d�'�4����K����[��d1��*���
�:�%�d����������9��d��U���u�u�u�u�w�4�(���;����lW��1����m�u�h�<���5�������9��h_�B���n�u�u�u�w�}�W���Yӏ��K5��N!��*���0�
�d�l�k�}� ���,����G9��Q��E���%�n�u�u�w�}�W���Y����V
��Z�*���
�d�a�i�w�8�(���H����lW�� 1��N���u�u�u�u�w�}�Wϭ�����R��R	��D���i�u�0�
�:�l�(���H����CT��N��U���u�u�u�u�$�1����L����lT��N�U���
�8�d�
�"�l�Oց�K���F�N��U���u�&�9�!�'�k����K����[��R����
� �d�l��o�}���Y���F�N�����!�%�b�'�0�o�B���Dӕ��l��Y�� ��e�
�g�_�w�}�W���Y���F��[1�����'�2�g�`�w�`��������l ��_�*��_�u�u�u�w�}�W���Y����G��1����c�u�h�&�;�)��������U��UךU���u�u�u�u�w�}�����ד�V��V�I���0�
�8�d�1��Oځ�K���F�N��U���u�&�9�!�'�����I���F��[1��؊� �m�d�%�l�}�W���Y���F���*���f�'�2�g�n�}�Jϭ����� 9��hV�*��_�u�u�u�w�}�W���Y����G��h��*��g�i�u�0��0�C���&����CT��N��U���u�u�u�u�$�1����&����V��R�����!�%�
� �o�n���Y���F�N��U���0�
�8�m�%�:�E��Y����V
��Z�����b�
�g�_�w�}�W���Y���F��[1�����2�g�a�u�j�.����	����S��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����%�!�;�%�g�4�G�������C9��Y�����6�d�h�4��4�(�������C��D��*���
�|�4�1��-��������lV������1�
� �m�b�-�^�������F�N��U���u�u�<�
�>���������9��E��G��u�h�<�
�>���������9��Q��G���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�0�
�'�)����I����F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����&�2�
�&��t����Q����\��h��*���u�%�'�2�'�.��������WW��R	��E���%�e�<�d�~�}����Y���F�N��U���
�
� �3�%�l�(�������F���*���3�'�d�
�c�/���J��ƹF�N��U���u�u�
�
�"�;���&����T9��N�U���
� �3�'�f��C���&����l��=N��U���u�u�u�u�w��(�������9��h��*��u�h�%�a�5�;����M����A��\�N���u�u�u�u�w�}�WϮ�M����U��Z��C���2�b�a�i�w��(�������9��h��*��g�_�u�u�w�}�W���Y�Ƽ�9��Q��*���g�'�2�c�a�a�W���&����V��1�����g�e�n�u�w�}�W���Y�����h�����d�
�
�0��k�W��	�ғ�F ��E1�*Ҋ�0�
�g�g�]�}�W���Y���F�G1�����0�
�a�l�%�:�A��E�Ƽ�9��Q��*���d�
�0�
�e�j�}���Y���F�N�����7�3�0�
�c�/���I���C9��U�����a�d�'�2�e�m�L���Y���F�N��U���
� �3�'�f��(���&����[��hZ�� ���'�d�
�d�%�:�E��B���F�N��U���u�
�
� �1�/�Fځ�M����lQ��R�����7�3�0�
�b�o�(���H����CU��N��U���u�u�u�u�'�i��������lW��E��B��i�u�
�
�"�;���&�ד�F9��^��F�ߊu�u�u�u�w�}�W���&ǹ��U ��h_��G���2�c�l�i�w��(�������9��E��G��n�u�u�u�w�}�W���YӖ��l��Q��Dߊ�
�0�
�b�w�`��������A9��hV�����g�g�_�u�w�}�W���Y���C9��U�����`�l�'�2�`�l�K���&ǹ��U ��h_��Dي�0�
�g�b�]�}�W���Y���F�G1�����0�
�`�'�0�k�D��Y����Q��R��@���'�2�g�a�l�}�W���Y���F���*���3�'�d�
��8�(��Y����lR��B����
�d�3�
�`�m���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������Z��h��*���|�4�1�}�/�)����&����V��S�����;�!�9�d�g�}��������]��[����h�4�
�<��.����&����@��h��*���|�!�0�_�w�}�W���Y���F��1�����
�a�d�
�2��E��E�Ƽ�9��Q��*���d�
� �d�`��D�ԜY���F�N��Uʥ�a�7�3�0��i�F�������F���*���3�'�d�
��(�F��&����F�N��U���u�u�%�a�5�;����M�ғ�V��^�I���
�
� �3�%�l�(ہ�����9��d��U���u�u�u�u�w�-�C�������R��h��*��g�i�u�
��(����Hǹ��U��Z����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�8�����ד�V��]�Hʴ�
�:�&�
�!��^Ͽ��έ�l��D�����
�u�u�%�$�:����&����CV��C	�����d�u�;�u�6�����&����P9��
N��*���
�%�!�;�'�m���P�Ƹ�VǻN��U���u�u�u�u����������W��R	��G��i�u�
�
�"�;���&�ד�F9��[��F�ߊu�u�u�u�w�}�W���&ǹ��U ��h_��G݊�0�
�g�b�k�}�(ہ�����lW��Y�� ��a�
�f�_�w�}�W���Y���F��1�����
�a�f�
�2��E��E�Ƽ�9��Q��*���f�
� �d�n��D�ԜY���F�N��Uʥ�a�7�3�0��i�Cށ����� Q�
N��A���3�0�
�a�c����Mƹ��l�N��U���u�u�u�%�c�?����&�ӓ� 9��P1�@���h�%�a�7�1�8�(���H����lW��1��N���u�u�u�u�w�}�WϮ�M����U��[��*���
�g�g�i�w��(�������9��Q��@���%�n�u�u�w�}�W���Y����lR��B����
�
�0�
�e�j�K���&ǹ��U ��h_��A���
�`�c�%�l�}�W���Y���F���*���3�'�d�
��8�(��K���C9��U�����`�m�3�
�b�j���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ڊ�!�g�3�8�d�}��������]��[����h�4�
�0��-����	�֓�GV�V ��]���!�:�1�
�2��G��DӇ��P	��C1��D��|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����<�0�
�%��)�^Ͽ��Ω�Z��Y
�����g�f�u�u�'�>�����ד�F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����&�2�
�&��t�^�����ƹF�N��U���u�u�0�
�d�}�JϹ�	����U��G_�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������%�<�0�
�'��������V��T��D���2�g�f�u�w�-��������lV�V ��]���6�;�!�9�0�>�F������T9��R��!���e�&�2�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۃ��G��S_�����e�b�h�4��2����¹����F��*���&�
�:�<��}�W���
����@��d:��ڊ�!�e�3�8�f�}��������]��[����h�4�
�0��-����	�֓�GW�G�����u�u�u�u�w�}�W�������W�
N�����
�g�
�g�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�!�0�9�%�W�������C9��h��\ʺ�u�=�u�!�#�}�������l�N��*���3�8�4�&�0�����CӖ��P��F��*���3�8�u�%�4�q��������Z��h��*���y�4�
�0��-����	�֓�GW�V�����1�
�b�y�2�4����H����R��G\����<�
�&�$���߁��ד�@��d��Uʷ�2�;�u�u�w�}����Y����`9��ZN�����u�u�u�u�w�5�Ͽ�&����GW��D��U��_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\��G1�����1�c�c�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����CV��C	�����d�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��E���8�d�h�u�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����V��G�����e�<�e�u�9�}��������]��[��E��0�<�6�;�f�;�(��&����� ��]´�
�:�&�
�8�4�(���Y����V��G�����e�<�d�|�~�t����s���F�N��U���u�u�4�
��;���Y����g9��1��ۊ�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�m�3�8�b�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��G�����
�&�
�u�i�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1�����
�%�
�!�~�<����	����@��X	��*���u�%�&�2�4�8�(���	�֓�G��Q��G���;�u�:�}�6�����&����P9��
N��*���
�%�!�;�'�m���P�����Yd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���%�e�&�2��.�(��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�O�������F�N��U���u�u�0�1�>�f�W���Y���F��_������%�e�&�0�����Y���F�N��U���u�u�4�
��;���Y����g9��1��ي�&�
�n�u�w�}�W���Yӑ��]F��h=�����&�2�
�&��}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����@��h��*��u�u�u�u�w�}� ���Y����g9��1�����h�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�;���s���F�N�����u�!�0�&�j�}�}���Y���F�N������3�8�i�w��/���[���F�N��ʶ�&�n�u�u�2�9��������9F�C����:�0�4�&�0�}����
���l�N��*���0�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���&����OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���A����lS�N�����u�u�u�u�w�}�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�1�;�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�4����
������T��[���_�u�u�%�>�1�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�_�u�w�8��ԜY���F��F�����4�
�:�&��2����Y�ƭ�l��E��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�%�<�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����0�1�u�&�>�3�������KǻN�����4�,�4�&�0�����CӖ��P�������4�
�<�
�$�,�$���˹��^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����u�u�u�u�w�}�WϿ�&����JF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�2�9�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�A���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�f�i�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ڊ�
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����H�ƭ�@�������{�x�_�u�w�-��������U��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�d�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�o�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(ց�	����l�N�����u�u�u�u�w�}�W�������T9��S1�G��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�I�ߓ�C9��SG����u�;�u�'�4�.�L�ԶY���F��h��*���
�f�u�&�>�3�������KǻN�����2�7�1�d�f�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�e�d��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����U��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m�F߁�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��D��4�&�2�u�%�>���T���F��h��*���
�a�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1�U���
�d�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����H���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�f�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��W�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��D؊�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��C���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�e�d�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��V�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lV��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�o�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���K�ƭ�@�������{�x�_�u�w�-��������T��V�����'�6�o�%�8�8�ǿ�&����P��h=�����&�2�
�&��q��������l ��Z�����u�u�7�2�9�}�W���Y���F������7�1�d�g�w�`�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���	ù��TV��D��\ʴ�1�;�!�}�'�>�����ד�[��O�����
� �m�`�'�t�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Y�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lV��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�`�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���OӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ù��l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�b�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��[�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��l�W�������A	��D�X�ߊu�u�%�&�0�?���N����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��D���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�g�u�&�>�3�������KǻN�����2�7�1�g��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��E����C9��h��]���:�;�:�e�w�}��������EW��UךU���;�u�'�6�$�f�}���Y���R��^	�����g�u�&�<�9�-����
���9F������7�1�g�c�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�b�d�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
����������F�R �����0�&�_�_�w�}�ZϿ�&����Q��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*؊�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��D���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�b�g�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��V�����u�u�7�2�9�}�W���Y���F������7�1�g�a�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��hY��*���#�1�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��B���
������T��[���_�u�u�%�$�:����K�Փ�@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q����M����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����9��h��\��u�u�0�1�'�2����s���F������7�1�g�g�6�.��������@H�d��Uʴ�
�<�
�1��k�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
���������F��P��U���u�u�u�u�w�}��������W9��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�@�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�g�d�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b�c�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����K���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Mڊ�&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��hY��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��e�W��Q����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����b�4�
�9�~�f�W�������A	��D����u�x�u�%�$�:����K����@��YN�����&�u�x�u�w�<�(���&����^��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�g�l�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������hV�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��d�W�������A	��D�X�ߊu�u�%�&�0�?���A����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�@�������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��L���h�}�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O��Y
�����:�&�
�:�>��W���&Ĺ��R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�f�b�4�$�:�W�������K��N�����<�
�1�
�g���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�g�<�(���P�����^ ךU���u�u�u�u�w�}��������lU��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(�������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��u�&�<�;�'�2����Y��ƹF��G1�����1�f�c�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�b�d�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�b�f���������F�R �����0�&�_�_�w�}�ZϿ�&����Q��\����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�D��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�g�4��1�^��Y����]��E����_�u�u�x�w�-�������� R��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��]�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��]�����1�_�u�u�2�4�}���Y���F�N�����<�
�1�
�d�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��B��
�%�#�1�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������U��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�ѓ�9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�f�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h_�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�EϿ�
����C��R��U���u�u�4�
�>�����L����@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(؁�L����E
��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����S��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�n�F���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�n�m������ƹF��R	�����u�u�u�u�w�}�W���
����W��_��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����e�4�&�2�w�/����W���F�V�����1�
�b�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�l�f�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W�� W�����;�%�:�0�$�}�Z���YӇ��@��U
��F���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��G���
�9�|�u�w�?����Y���F�N��U���%�&�2�7�3�n�N��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lU��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��lU��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����9�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�@Ͽ�
����C��R��U���u�u�4�
�>�����@Ĺ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ց�&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��F��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ�l��A��\�ߊu�u�;�u�%�>���s���K�V�����1�
�e�u�$�4�Ϯ�����F�=N��U���&�2�7�1�c�k��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�l�b�<�(���P�����^ ךU���u�u�u�u�w�}��������lR��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(ځ�	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��A���&�<�;�%�8�8����T�����D�����a�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ڊ�
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��E���R��X ��*���<�
�u�u���(������R��Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��[�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����l_��h�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�d�w�`�_���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1��C���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&Ĺ��l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����a�i�u�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�N�����%�6�;�!�;�:���DӖ��lQ��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�f�w�.����	����@�CךU���%�&�2�7�3�i�D���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�n�e������ƹF��R	�����u�u�u�u�w�}�W���
����W��]��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����g�4�&�2�w�/����W���F�V�����1�
�a�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&����[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�l�n�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��_�����;�%�:�0�$�}�Z���YӇ��@��U
��A���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1��Dڊ�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��B���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�l�d�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��^�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����l_��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�g�a�Wǰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�4�1�}�'�>��������lW���*���4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ʹ��l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�c�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��\�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��j�W�������A	��D�X�ߊu�u�%�&�0�?���A����Z��G��U���'�6�&�}�'�.����Y����Z��D��&���!�
�&�
�{�-�N��&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��A��i�u�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ߓ� 9��h��\��u�u�0�1�'�2����s���F������7�1�a�b�6�.��������@H�d��Uʴ�
�<�
�1��e�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��i������ƹF��R	�����u�u�u�u�w�}�W���
����W��Y��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ց�M����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����l�u�&�<�9�-����
���9F������7�1�a�c�6�.���������T��]���&�4�!�u�'�.��������l��h��*���%�l�d�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�n�l�(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�U���<�;�%�:�2�.�W��Y����C9��P1�����
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*ۊ�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��G��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lS��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�d�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lS��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�%�4�3����H�����t=�����u�:�;�:�c�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lS��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�f�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����_��D�����:�u�u�'�4�.�_���
����F��h��*���$��
�!��.�(��	�֓�l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�l�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lV��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�`�}����Ӗ��P��N����u�%�&�2�5�9�A�������]9��X��U���6�&�}�%�$�<����&ù��R��[
�����2�u�
�
��-��������TJ��h^��*���#�1�<�
�>�q����J����E
��^ �����%�e�a�4��1�(���
���C9��1��*���
�;�&�2�w��(ف�	����l��D��U���
�
�%�#�3�4�(���UӖ��l^��G1�����
�<�y�%�g�d��������l��N��E��
�%�#�1�>����	�֓�9��h��*���&�2�u�
��o��������l��N��E��
�%�#�1�>����	�֓�9��h��*���&�2�u�
��h��������l��N��B���4�
�9�
�9�.����&Ĺ��R��[
�����2�u�
�
��-��������TJ��hY��*���#�1�<�
�>�q����M����E
��^ �����%�b�`�4��1�(���
���C9��1��*���
�;�&�2�w��(؁�	����l��D��U���
�
�%�#�3�4�(���UӖ��l_��G1�����
�<�y�%�`�l�(�������]9��PB��*݊�d�4�
�9��3����Y����T��G1�����
�<�y�%�`�l�(�������]9��PB��*݊�a�4�
�9��3����Y����S��G1�����
�<�y�%�n�m��������l��N��L���4�
�9�
�9�.����&ʹ��R��[
�����2�u�
�
��-��������TJ��hW��*���#�1�<�
�>�q����L����E
��^ �����%�l�c�4��1�(���
���C9�� 1��*���
�;�&�2�w��(ׁ�	����l��D��U���
�
�%�#�3�4�(���UӖ��lW��V�����;�&�2�u���F���&����Z��^	����d�
�%�#�3�4�(���UӖ��lW��V�����;�&�2�u���C���&����Z��^	����d�
�%�#�3�4�(���P�����^ ךU���u�u�u�u�w�}��������lP��R��]¥�l�e�4�
�;���������C9��Y�����6�e�u�'���(ށ�	����l��D��Hʴ�
�:�&�
�8�4�(�������l_��h�����<�
�<�u�w�-��������Z��N��U¥�l�f�4�
�;���������C9��Y�����6�e�u�'���(ہ�	����l��D��Hʴ�
�:�&�
�8�4�(�������l_��h�����<�
�<�u�w�-��������Z��N��U¥�l�c�4�
�;���������C9��Y�����6�e�u�'���(؁�	����l��D��Hʴ�
�:�&�
�8�4�(�������l_��h�����<�
�<�u�w�-��������Z��N��U¥�l�l�4�
�;���������C9��Y�����6�e�u�'���(�������W9��h��U���%�6�;�!�;�:���Y���C9��_�����1�<�
�<�w�}��������\��h^�����%�l�d�
�'�+����&����F��h�����:�<�
�|�8�}����H����l��h�����h�4�
�:�$�����&����AF��hW��A���
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�b�<�(���&����Z������!�9�2�6�g�}����&Ĺ��R��[
�����2�h�4�
�8�.�(�������	����*ۊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�b�e�<�(���&����Z������!�9�2�6�g�}����&Ĺ��R��[
�����2�h�4�
�8�.�(�������	����*ފ�%�#�1�<��4�W���	����@��X	��*���:�u�%�b�b�<�(���&����Z������!�9�2�6�g�}����&Ĺ��R��[
�����2�h�4�
�8�.�(�������	����*݊�%�#�1�<��4�W���	����@��X	��*���:�u�%�b�o�<�(���&����Z������!�9�2�6�g�}����&Ĺ��R��[
�����2�h�4�
�8�.�(�������	����*���4�
�9�
�9�.�������]��[����u�'�}�
��l��������l��S�����;�!�9�2�4�m�W���Q����T��G1�����
�<�u�u�'�>��������lV�X�����d�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�j�Fہ�	����l��D��Hʴ�
�:�&�
�8�4�(�������lQ��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G�������W9��h��U���%�6�;�!�;�:���Y���C9��1��*���
�;�&�2�j�<�(���
����T��G�����
�
�
�%�!�9�������R��X ��*���<�
�|�:�w�-�G��&����_��Y1����4�
�:�&��2����PӉ����h_�����9�
�;�&�0�`��������_	��T1�U���}�
�
�g�6���������[��G1�����9�2�6�e�w�/�_���&�Փ�C9��S1��*���u�u�%�6�9�)�������\�G1��Dފ�%�#�1�<��4�W���	����@��X	��*���:�u�%�e�f���������@��
N��*���&�
�:�<��t��������R��
N��*���&�
�:�<��t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������T9��R��!���d�3�8�e�w�-��������P�N�����;�u�u�u�w�}�W���YӇ��@��U
��C��i�u�}�%�4�3��������[��G1�����0�
��&�f�;���Y����]	��V�����1�
�b�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y���� 9��h��\��u�u�0�1�'�2����s���F������7�1�b�u�$�4�Ϯ�����F�=N��U���&�2�7�1�`���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����Q�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���(������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�Gʴ�&�2�u�'�4�.�Y��s���R��^	�����a�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�c�}�J���	����@��A_��U���%��
�&��}�������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�U���<�;�%�:�2�.�W��Y����C9��P1����
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*ߊ�%�#�1�_�w�}����s���F�N��U���4�
�<�
�3��A��Yۈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�4�3�u��������\��h_��U���
�
�%�#�3�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������l_��h�����%�:�u�u�%�>��������]��E��G��y�4�
�<��.����&����@��h��*���4�
�0�
�'�)����I����l�N�����u�u�u�u�w�}�W�������T9��S1�G��u�}�-�!�8�9�(���&����[��G1�����9�d�e�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����l ��h_�����}�%�6�;�#�1����H����C9��P1�����
�%�
�!�~�f�W�������A	��D����u�x�u�%�$�:����@����@��YN�����&�u�x�u�w�<�(���&����
W��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��L��i�u�4�
�8�.�(���&���R��d1�����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����@�ƭ�@�������{�x�_�u�w�-��������9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&ù��R��[
��U���7�2�;�u�w�}�W���Y�����D�����l�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��V�����n�u�u�0�3�-����
��ƓF�C�����2�6�0�
��-�G���ù��^9��V�����'�6�&�{�z�W�W���	����l��F1��*���
�!�e�3�:�l��������\������}�%�&�2�5�9�B��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��E���8�d�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���%�e�&�2��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ڊ�!�d�3�8�e�<����Y����V��C�U���4�
�<�
�$�,�$���	ù��TW��D��*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�m�g�u�?�3�}���Y���F�V�����&�$��
�'���������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l��1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���&����l ��h]�����;�%�:�0�$�}�Z���YӇ��@��T��*���%�e�&�2��.�(܁�
����l��TN����0�&�4�
�>�����M��ƹF��R	�����u�u�u�3��-��������V�C��U���u�u�u�u�w�<�(���&����l5��G�����
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�%�
�#�o����J���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���e�&�2�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l��1�����4�&�2�
�%�>�MϮ�������D�����`�c�_�u�w�8��ԜY���F��F��*���
�1�
�`�~�)����Y���F�N�����2�6�0�
��-�G�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������C��D��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ד�@�������%�:�0�&�w�p�W�������T9��R��!���d�3�8�e�6�.���������T��]���&�2�7�1�e�t�W�������9F�N��U���}�%�&�2�5�9�E�������9F�N��U���u�%�&�2�4�8�(���
�ד�@��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��M���8�`�4�&�0�����CӖ��P�������7�1�l�b�]�}�W������F�N��U´�
�<�
�1��l�^Ϫ���ƹF�N��U���%�&�2�6�2��#���A����lS�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����G^��D��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��O�����
� �m�`�'�}�J���[ӑ��]F��{1��*���
�:�%�`�'�4����K����[��G1�����9�`�d�|�2�.�W��B��� ��[�����:�%�d�
��5�(���H����CU�
NךU���u�u�
�
��3����������h��F���
�l�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�d��(�F��&����F�Q=�����'��:�
�c�l��������V��N�U���u�u�u�%�n�l�����ƻ�V�D�����l�3�
�d�d�-�_���D����F��D��U���u�u�&�9�#�-�B���&����l��=N��U���u��;�1��8��������
_��N�U���
�:�<�
�2�)�Ǭ�
����@��R
��"��� �,� �
��8�(��@����O��=N��U���u��;�1��8���&����lW��1��U��&�1�9�2�4�+����Q����I��^	��¼�
����#�l�(ށ�����T�\��N�ߠu�u�x�u�%����@����R��P �����&�{�x�_�w�}��������l��V�����'�6�o�%�8�8�ǿ�&����C��R ��ڊ�!�y�4�
�>�����*����9��P]�����y�4�
�<��.����&����@��h��*���4�
�0�
�'�)����I����F��h��3����:�
�a�g�-��������J��d1��*���
�:�%�d����������Q�N�����;�u�u�u�w�4�W�������]��[����h�4�
�<��.����&����@��h��*���4�1�}�%�4�3��������[��G1�����<�0�
�%��)�^�������9F�N��U���u�'�
� �o�d����DӀ��_��X�����d�
�
�=��8�(��N���F�N�����}�}�%�6�9�)���������E�����0�
�%�
�#�t����Q����\��h�����u�u�%�&�0�>����-����l��1����|�u�=�;�]�}�W���Y���T��Q��Gӊ�e�i�u��;���������9��G�����g�e�n�u�w�}�Wϻ�
��ƹF�N��U���'�
� �m�n�-�W��[����k>��o6��-���������/���[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�f�
�2�<����Y����V��C�U���2�%�3�
�d�����
����C��T�����&�}�%�6�{�<�(���&����l5��G�����
�&�
�y�6�����
����g9��1��ي�&�
�y�4��4�(�������C��D��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R��F��*���&�
�:�<��}�W���
����@��d:��ڊ�!�g�3�8�d�}����	����@��X	��*���u�%�&�2�4�8�(���	�֓�G��Q��A���'�}�%�6�9�)���������D�����
��%�e�$�:�(���&���F��R ��U���u�u�u�u�0�-����J����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�'�
�"�e�D���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z�������l^��h����2�u�'�6�$�s�Z�ԜY�ƫ�C9��hV�*���4�&�2�
�%�>�MϮ�������D�����
��%�e�$�:�(���&����C9��P1�����
�%�
�!�{�;�(�������^9��Q��G���%�y�4�
�>�����*����9��P_�����y�3�
�:�2�)����M����F9��]��D�ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�6�����	����l��h��\���=�;�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��h��G���8�f�|�!�2�}�W���Y���F�N����� �m�f�%�w�`��������V��Z��*���d�e�
�d�]�}�W���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���
�!�d�3�:�o�^Ϫ���ƹF�N��U���u�u�'�
�"�e�D���Y����`9��S�����f�3�
�g�n�-�L���Y���F����ߊu�u�u�u�w�}�W�������l^��h�I���������/���!����k>��o6��-���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���0�_�u�u�w�}�W�������l^��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�>���������C9��1�E���3�
�e�d�'�}�J�������l^��h����%�6�;�!�;�i�F��Y����9��h(��*���%�`�d�d�1��E���	�����h�����0�!�'� �$�:����	����@��A[��\��� �&�2�0����������\��h��*���m�g�%�|�l�W�W���Tӏ��_��X�����`�%�<�3��o�(������]F��X�����x�u�u�<��4�1���5����9��^1��*��
�a�4�&�0�����CӖ��P�������:�
�:�%�b�/���A�Ʃ�Z��Y
�����g�f�y�4��4�(�������C��D��*���
�y�4�
�2���������l��N��*����'��:���(ށ�����Q�N�����;�u�u�u�w�4�W�������\��h��*��b�h�4�
�8�.�(���&����]�V�����
�:�<�
�w�}��������B9��h��*���e�3�8�d�w�3�Wǿ�&����G9��P��D��4�
�0�
�'�)����I����O�C��U���u�u�u�u�w�4�(���?����\	��1�����
�g�
�a�k�}�;���&����	��h[��*ۊ�0�
�d�b�]�}�W���Y����l�N��U���u�<�
�<��/�;���&ƹ��Z9��hV�*��i�u��9��2�(���	�ӓ�V��V�U���u�u�0�1�>�f�}���Y����C��R�����u�<�
������&¹��lW�� 1��U��&�1�9�2�4�+����Q����T�� ��&���e�3�
�d�d�-�^������]��Y����
� �d�f��n�^�ԜY�ƥ�l��u�����3�
�e�`�'�}�Jϭ�����Z��R�� �&�2�0�}�2��ف�����l��C�����;�1�;�"�2�l�(���H����CU�d��Uʻ�"�0�d�
�"�d�@���Y���F�N�����g�<�
�<�w�5��������C9��hV�*��e�u�u�d�~�8����Y���F��hY��A���
�<�n�u�w�3� ���H¹��l_��h�I���u�u�u�u�9�*��������
9�������'�6�;�
�"�d�D���Q���A��N�����u�u�u�u�9�*��������9��d��Uʻ�"�0�d�
�"�l�Gށ�J���9F�N��U����9�
� �n�l�������\��X ��*���l�b�%�}�~�`�P���Y����l�N��Uʻ�"�0�d�
�"�d�@���B�����d��F���
�e�l�%�w�`�}���Y���]��R�*���l�f�%�u�?�3�_�������l ��Z�����|�h�r�r�w�1��ԜY���F��@=��D؊� �d�e�
�d�W�W�������R��B1�Dӊ�f�i�u�u�w�}�WϮ�I�ד�]9��PN�����&�9�!�%�n�;�(��J����O�I�\ʰ�&�u�u�u�w�}����H����l��d��Uʻ�"�0�d�
�"�l�Dށ�J���9F�N��U���
�d�<�
�>�}����Q����G�� 1��*��d�%�}�|�j�z�P������F�N�����l�<�
�<�l�}�Wϰ�����9��h_�F���u�h�_�u�w�}�W���&Ĺ��l�������0�
�8�d��(�F��&���F�_��U���0�_�u�u�w�}�(߁�&����Z��N�����0�d�
� �f�h�(��E��ƹF�N��*ڊ�
�;�&�2� �8�Wǭ�����U��B1�B݊�g�e�u�u�f�t����Y���F���*���<�
�<�n�w�}��������U��X�����h�_�u�u�w�}�����ғ�F9��W��Fʢ�0�u�:�
�8�9�(���H����CT�N��R��u�9�0�_�w�}�W�������S��B1�Fۊ�f�_�u�u�2���������S��N�U���u�u�u�;� �8�Fف����� 9�������'�6�;�a�1��F���	����[�I�����u�u�u�u�w�3� ���HĹ��lW��1��N���u�;�"�0�f�;�(��&���FǻN��U���
�
�e�<��4�W����ο�_9��GV�� ��l�%�}�|�j�z�P������F�N�����m�<�
�<�l�}�Wϰ�����9��h_�F���u�h�_�u�w�}�W���*����l ��_�*��"�0�u�:��2�ځ�����
9��^��H��r�u�9�0�]�}�W���Y����V
��h��D��
�f�_�u�w�8�$���H����W��h�I���u�u�u�u�'�j�F���&����D��F�����%�l�3�
�f�n����P���A�R��U���u�u�u�%�`�l�(���
����F�Y����
� �d�l��n�K���Y���F��hY��D���
�<�u�=�9�u��������U��^�����|�h�r�r�w�1��ԜY���F�� 1�����<�n�u�u�9�*���&����V��G]��H�ߊu�u�u�u���(���
����[����*���d�
� �d�o��E��Y���O��[�����u�u�u�
���������F��@=��Gފ� �d�e�
�d�a�W���Y�����h]�����2�"�0�u�$�1����J����V��h�E���u�d�|�0�$�}�W���Y����lQ��1��*���n�u�u�;� �8�Eځ�����9��R�����u�u�u�0��1�F���&����l��@��Uº�
�:�1�
�"�l�Eځ�K���F�G�����_�u�u�u�w�8�$���K����W��h����u�0��9�a�;�(��J����[�N��U���;�"�0�g��(�F��&����[�������a�3�
�d�n�-�_���D����F��D��U���u�u�;�"�2�o�(���H����CU��N�����0�g�
� �f�n�(��E��ƹF�N�����9�`�3�
�e�h�������\��X ��*���d�c�
�g�g�}�W��PӃ��VFǻN��U���0��9�c�1��E���	��ƹF��R��؊� �l�d�%�w�`�}���Y���C9��1��*���u�=�;�}�2���������9��^��H��r�u�9�0�]�}�W���Y����9��h��N���u�;�"�0�d�;�(��&���FǻN��U���
�
�
�;�$�:� ���Yە��l��h��M���%�}�|�h�p�z�W������F�N��E��
�;�&�2�]�}�W���*����U��W��F��u�u�u�u�w�3� ���&����
Q��N�����:�
�:�1�1��G܁�K���F�G�����_�u�u�u�w�8�$���&����_��UךU���0��9�
�"�d�D���Y���F�N�����0�g�3�
�e��Dϩ�����A9��Y
�����g�
�g�e�w�}�F�������9F�N��U����9�
� �n�n���Y����V��[X�� ��d�%�u�h�]�}�W���Y����V
��Q��Fӊ�f�"�0�u�8�����&����Q��F�U���d�|�0�&�w�}�W���Yӈ��`��h��L���%�n�u�u�9�*��������
9��R�����u�u�u�
������ӑ��]F��R�����3�
�l�
�e�m�W���H����_��=N��U���u�
�
�g�>����Y����V��[V�� ��`�%�u�h�]�}�W���Y����V��Y1��ʢ�0�u�&�9�#�-�(���A�ߓ�N��S��D���0�&�u�u�w�}�WϮ�N�ޓ�]9��PUךU���0��9�
�"�d�F���Y���F�N�����c�<�
�<�w�5��������CR��B1�B���}�|�h�r�p�}����s���F�G1��A���
�<�n�u�w�3� ���&����
Q��N�U���u�u�u�%�g�m�����ƻ�V�D�����
� �m�d�'�u�^��^���V
��d��U���u�%�e�d��3����s���\��X ��*���l�`�%�u�j�u�����ޓ�F9��1��U���&�9�!�%��(�O���	����F�X�����
� �l�b�'�}�J�������CR��B1�B���u�'�&�9�#�-�(���A�ד�O��N�����:�1�
� �n�j����D�Σ�l��S1��*��
�g�:�u�%�>��������9��UךU���'�6�;�a�1��F���	���N��[1�����3�
�e�l�'�}�ϭ�����R��B1�Mي�g�n�u�u�8�����&����P��G\��H���'�6�;�m�1��F���	�ƣ�	��T��L���
�d�b�%�~�W�W�������W^��B1�Gߊ�g�i�u�&�;�)��������U��N��U���
�8�d�
�"�l�G؁�K��ƹF��E1�����3�
�d�b�'�}�J�������CW��Q��D���%�u�'�&�;�)��������
S��G�U���:�
�:�1�1��G܁�K�����h��F���
�l�
�g�8�}�����ד�F9��1��\�ߠu�u�x�u���(�������]9��PN�����u�'�6�&�y�p�}���Y����9��h��*���&�2�4�&�0�����CӖ��P����*ڊ�%�#�1�u���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�e�e�6�����Y����l�N��U���u�%�e�e�6���������Z�G1��E���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�%�!�9���������h^�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lV��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�&�<�;�'�2�W�������@N��1�U���
�
�'�2�w��(߁�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�;�$�:�K���&ù��9F�N��U���0�_�u�u�w�}�W���&ù��Z��^	��Hʥ�e�e�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lV��1��*���
�;�&�2�6�.��������@H�d��Uʥ�e�d�
�%�!�9��������@��h����%�:�0�&�'�m�F߁�	����F��1�*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��h�����|�!�0�u�w�}�W���Y����lV��1��*���
�;�&�2�k�}�(߁�I����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��h�����<�
�<�u�j�-�G��&����_��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���G���&����R��P �����&�{�x�_�w�}�(߁�I����@��V�����'�6�o�%�8�8�Ǯ�I������h_�����y�%�e�d��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���4�
�9�|�w�5��ԜY���F�N��E��
�;�&�2�k�}�(߁�I���F�N�����u�u�u�u�w�}����Hù��l��R�����d�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�d�4�
�;���������Z��G��U���'�6�&�}���F���&������h_�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lW��V�����u�=�;�_�w�}�W���Y�Ƽ�9��h�����<�
�<�u�j�-�G��&����_��N��U���0�&�u�u�w�}�W���YӖ��lW��V�����;�&�2�i�w��(�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g�l�(���
����@��YN�����&�u�x�u�w�-�G��&����Z��D�����:�u�u�'�4�.�_���&���C9��_�����u�
�
�d�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��Dۊ�%�#�1�|�#�8�W���Y���F���*���<�
�<�u�j�-�G��B���F����ߊu�u�u�u�w�}�(߁�H����@��S��*ڊ�d�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lW��V�����;�&�2�4�$�:�W�������K��N�����d�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�g�l�(������C9��\�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����T��G1�����!�0�u�u�w�}�W���YӖ��lW��V�����;�&�2�i�w��(�������W]ǻN��U���9�0�_�u�w�}�W���Y����T��G1�����
�<�u�h�'�m�F݁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��o�����ƭ�@�������{�x�_�u�w��(�������T9��D��*���6�o�%�:�2�.����H����lV��1�����%�e�d�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h^��G���
�9�|�u�?�3�}���Y���F�G1��D؊�;�&�2�i�w��(��s���F�R��U���u�u�u�u�w�-�G��&����Z�
N��E��
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����U��G1�����
�<�u�&�>�3�������KǻN��*ڊ�f�4�
�9��3��������]9��X��U���6�&�}�
��n��������lV��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�֓� 9��h��\���=�;�_�u�w�}�W���Y����U��G1�����
�<�u�h�'�m�F܁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�֓� 9��h��*���&�2�i�u���D���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e�f�����Ӈ��Z��G�����u�x�u�u�'�m�F܁�����l��^	�����u�u�'�6�$�u�(߁�J�Ƽ�9��h�����
�
�f�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�*���#�1�|�!�2�}�W���Y���F��h^��F���
�<�u�h�'�m�F��Y���F��[�����u�u�u�u�w��(�������TF���*���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�֓�9��h��*���&�2�4�&�0�}����
���l�N��E��
�%�#�1�>�����
����l��TN����0�&�%�e�f������Ƽ�9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��l��A��\ʡ�0�u�u�u�w�}�W���	�֓�9��h��*���&�2�i�u���C���&����9F�N��U���0�_�u�u�w�}�W���&ù��l��A�����<�u�h�%�g�l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�c�4�(���Y����T��E�����x�_�u�u���C���&����R��P �����o�%�:�0�$�-�G��UӖ��lW��G��Yʥ�e�d�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h_�����9�|�u�=�9�W�W���Y���F��1�*���&�2�i�u���C�ԜY���F��D��U���u�u�u�u�'�m�Fہ�����Z�G1��Dފ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��l��A�����<�u�&�<�9�-����
���9F���*���4�
�9�
�9�.����
����C��T�����&�}�
�
�b�<�(���UӖ��lW��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�I����R��[
��U���;�_�u�u�w�}�W���&ù��l��A�����<�u�h�%�g�l�(�������F�N�����u�u�u�u�w�}�WϮ�I����R��[
�����2�i�u�
��h��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�e�d��3��������]F��X�����x�u�u�%�g�l�(���
����@��Y1�����u�'�6�&���(��Y����S��E��U���
�`�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��[�����1�|�!�0�w�}�W���Y�����h_�����<�u�h�%�g�l�L���Y�����RNךU���u�u�u�u���B���&����[��h^��@���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�I�ד�C9��S1��*���u�&�<�;�'�2����Y��ƹF��h^��*���#�1�<�
�>���������PF��G�����%�e�d�4��1�[Ϯ�I�ד�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(ށ�	����O��_�����u�u�u�u�w��(ށ�	����l��D��I���
�
�
�%�!�9�}���Y���V
��d��U���u�u�u�%�g�l��������l��R�����d�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��D���
�<�u�&�>�3�������KǻN��*ڊ�
�;�&�2�6�.���������T��]���
�y�%�e�f�-���	�֓�l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g�l�������G��d��U���u�u�u�%�g�l���������h_�U���u�u�0�&�w�}�W���Y�����h_�����2�i�u�
������s���F�R ����_�u�u�;�w�/����B��ƹF�N��E���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e�e�<�(���&����Z��D�����:�u�u�'�4�.�_���&����l��N��E���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h\�����1�|�!�0�w�}�W���Y�����h\�����1�<�
�<�w�`����K����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��V�����;�&�2�i�w��(݁�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
������Ӈ��Z��G�����u�x�u�u�'�m�E���&����R��P �����o�%�:�0�$�-�G��Y����9��R	����g�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��^ �����h�%�e�g�]�}�W���Y����l�N��U���u�%�e�g�>�����DӖ��lT��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(�������]9��PN�����u�'�6�&�y�p�}���Y���� 9��h��*���&�2�4�&�0�����CӖ��P����*ي�%�#�1�u���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�e�f�6�����Y����l�N��U���u�%�e�f�6���������Z�G1��F���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�%�!�9���������h]�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lU��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�&�<�;�'�2�W�������@N��1�U���
�
�'�2�w��(܁�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�;�$�:�K���&ù��9F�N��U���0�_�u�u�w�}�W���&ù��Z��^	��Hʥ�e�f�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lV��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�g�i��������lV��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ù��R��[
��U���;�_�u�u�w�}�W���&ù��R��[
�����2�i�u�
���������F�N�����u�u�u�u�w�}����M����E
��^ �����h�%�e�a�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�e�a�<�
�>�}����Ӗ��P��N����u�
�
�
�9�.����
����C��T�����&�}�
�
�{�-�G���	������hZ�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����M����E
��N�����u�u�u�u�w�}����M����@��S��*ڊ�n�u�u�u�w�8����Y���F�N��*ڊ�
�;�&�2�k�}�(߁�&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�e�`�4��1�(���
����@��YN�����&�u�x�u�w�-�G�������W9��h��*���<�;�%�:�w�}����
�μ�9��V�����%�e�`�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ڊ�
�%�#�1�~�)����Y���F�N��*ڊ�
�%�#�1�>�����DӖ��lS��G1���ߊu�u�u�u�;�8�}���Y���F�G1��@���
�9�
�;�$�:�K���&ù��R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(߁�&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I�ӓ�]9��P1�����
�'�6�o�'�2����	�֓�F��1�����y�%�e�`�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��@���
�9�|�u�?�3�}���Y���F�G1��@���
�<�u�h�'�m�B�ԜY���F��D��U���u�u�u�u�'�m�B���&����[��h^��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&Ź��l��h�����4�&�2�u�%�>���T���F��1�����9�
�;�&�0�<����&����\��E�����
�
�
�%�!�9�W���&Ź��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�m�A���&����F��R ��U���u�u�u�u�'�m�A���&����Z��^	��Hʥ�e�c�4�
�;�f�W���Y����_��=N��U���u�u�u�
����������@��S��*ڊ�
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h^��*���&�2�4�&�0�}����
���l�N��E���<�
�<�
�$�4��������C��R�����c�u�
�
��/����&ù��R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
����������[��=N��U���u�u�u�
���������C9��UךU���u�u�9�0�]�}�W���Y���C9��1��*���u�h�%�e�a�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*݊�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��-��������T9��D��*���6�o�%�:�2�.����N����E
����*݊�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9�� 1��*���|�u�=�;�]�}�W���Y���C9�� 1��*���
�;�&�2�k�}�(߁�&����_��N��U���0�&�u�u�w�}�W���YӖ��lQ��G1�����
�<�u�h�'�m�@���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�e�`�4�(���Y����T��E�����x�_�u�u���(���
����@��Y1�����u�'�6�&���(��	�֓�l��PB��*ڊ�
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lQ��G1�����!�0�u�u�w�}�W���YӖ��lQ��Y1����u�
�
�n�w�}�W�������9F�N��U���u�
�
�
�9�.���Y����9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g�e��������l�������%�:�0�&�w�p�W���	�֓�l��A�����<�
�&�<�9�-����Y����V��G1��M���
�9�y�%�g�e��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�'�+��������9F�N��U���u�
�
�
�'�+����&����[��h^��*���#�1�_�u�w�}�W������F�N��Uʥ�e�m�4�
�;��������C9��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��h��U���<�;�%�:�2�.�W��Y����lV��h�����4�&�2�
�%�>�MϮ�������hV����m�%�0�y�'�m�O���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e�m�4�
�;�t�W������F�N��Uʥ�e�m�<�
�>�}�JϮ�I����F�N�����u�u�u�u�w�}�WϮ�I�ޓ�]9��PN�U���
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��V�����;�&�2�4�$�:�W�������K��N�����l�4�
�9��3��������]9��X��U���6�&�}�
�������Ƽ�9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�I�ߓ�C9��SG�����u�u�u�u�w�}�WϮ�I�ߓ�C9��S1��*���u�h�%�e�n�<�(���B���F����ߊu�u�u�u�w�}�(߁�&����_��Y1����u�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�;�&�0�<����Y����V��C�U���%�e�l�<��4�(�������A	��N�����&�%�e�l�w��(ց����C9��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(߁�&����_����ߊu�u�u�u�w�}�(߁�&����Z�
N��E��_�u�u�u�w�1��ԜY���F�N��E���<�
�<�u�j�-�G���	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*ފ�u�h�%�a�5�;����M����lP��dךU���x�%�a�e�6�����
������T��[���_�u�u�
����������Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=�����3�8�`�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)����Y���F�N��*ފ�
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h^�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����d�i�u�
��(����Hƹ��T9��UךU���
�
�e�i�w��(�������9��h��*��n�_�u�u�z�-�C��&����_��D��ʥ�:�0�&�u�z�}�WϮ�M����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�o�;���s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P����[��=N��U���u�u�u�
��m���������T�����2�6�d�_�w�}�W������F�N��U���%�a�d�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�i�F���DӖ��l��Q��Dߊ�a�'�2�b�d�W�W���T�Ƽ�9��h�����4�&�2�u�%�>���T���F��1�*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$���˹��^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ޓ�@��G�����u�u�u�u�w�}�WϮ�M����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w��(�������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����T�
N��A���3�0�
�g�$�/���O��ƹF�N��A��
�%�#�1�6�.��������@H�d��Uʥ�a�d�
�%�!�9��������\������}�%�6�y�6�����
����g9��1�����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��CV�����|�|�!�0�w�}�W���Y�����h_�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����T��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1��D���h�%�a�7�1�8�(���
����lQ��dךU���x�%�a�d��-��������]F��X�����x�u�u�%�c�l�(�������@��Y1�����u�'�6�&��-�������T9��R��!���m�3�8�`�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�t����Y���F�N��U���
�f�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1��Dي�%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�a�d�u�j�-�C�������R��h��*��n�_�u�u�z�-�C��&����_��D��ʥ�:�0�&�u�z�}�WϮ�M����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�o�;���s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P����[��=N��U���u�u�u�
��i���������T�����2�6�d�_�w�}�W������F�N��U���%�a�d�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�i�F���DӖ��l��Q��Dߊ�
�0�
�e�l�W�W���TӖ��lW��V�����&�<�;�%�8�8����T�����h_�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���A����lS�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9��G�����_�u�u�u�w�}�W���&�ӓ�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�i�Fځ�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lR��h�����4�&�2�u�%�>���T���F��1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���A����lS�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���˹��^9��G�����_�u�u�u�w�}�W���&¹��l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�M���F��1�����
�a�g�'�0�k�A�ԶY���F��1�����9�u�&�<�9�-����
���9F���*؊�%�#�1�4�$�:�(�������A	��D�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h[��\ʡ�0�u�u�u�w�}�W���	�ғ�l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�C�������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���� F���*���3�'�d�
��8�(��B���F���*ي�%�#�1�4�$�:�W�������K��N�����f�4�
�9��.����	����	F��X��´�
�0�u�%�$�:����&����G^��D��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��@���u�=�;�_�w�}�W���Y�Ƽ�9��V�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����lR��R�����7�3�0�
�c�h����O����9F�C����a�4�
�9�w�.����	����@�CךU���
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��1�����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��CV�����|�|�!�0�w�}�W���Y�����hZ�����1�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W���	�ғ�l��A��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��1�I���
�
� �3�%�l�(ځ�����]ǑN��X���
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�a�`�6�����
����l��TN����0�&�4�
�2�}��������B9��h��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��M���8�`�|�u�?�3�}���Y���F�G1��@���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��V�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*���h�%�a�7�1�8�(���@����lP��dךU���x�%�a�c�6�����
������T��[���_�u�u�
����������Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=�����3�8�`�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)����Y���F�N��*ފ�
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����hX�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����b�i�u�
��(����Hƹ��A�� ^����u�x�u�
������Ӈ��Z��G�����u�x�u�u�'�i�@���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�
�&�
�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�b�t�W������F�N��Uʥ�a�b�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1��B���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�u�h�'�i��������lW��E��B��_�u�u�x�w��(ׁ�	������^	�����0�&�u�x�w�}����A����E
��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�
�$��^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�m�1�0�B���Y����l�N��U���u�%�a�m�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����m�4�
�9�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�
�
�w�`��������A9��h_�����b�b�_�u�w�p�W���&ʹ��l�������%�:�0�&�w�p�W���	�ғ�l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�e����L���G��d��U���u�u�u�%�c�d���������T�����2�6�d�_�w�}�W������F�N��U���%�a�l�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u����������V��B1�Aӊ�f�i�u�u�w�}�WϹ�	����T��G\�����}�0�
�8�c�/���O����[�I�����u�u�u�u�w�-�C�������R��h��*��n�u�u�%�c�?����&�ғ�9��h_�C���u�h�_�u�w�}�W���&����V��1�����c�m�"�0�w�.����	����T9��\��\��r�r�u�9�2�W�W���Y�Ƽ�9��Q��*���d�
� �d�c��D�ԜY�Ƽ�9��Q��*���d�
� �d�a��D��Y���F���*���3�'�d�
��8�(��Y����N��[1�����2�g�a�}�~�`�P���Y����l�N��Uʥ�a�7�3�0��i�Fށ�����9��d��Uʥ�a�7�3�0��i�F܁�����9��R�����u�u�u�
��(����Hǹ��A��V����u�&�9�!�'�����I���F�_��U���0�_�u�u�w�}�(ہ�����lW��\�� ��c�
�f�_�w�}�(ہ�����lW��Y�� ��b�
�f�i�w�}�W���YӔ��l^�������0�
�8�c�%�:�E��Q���A��N�����u�u�u�u�'�i��������lW��E��B��_�u�u�
��(����Hǹ��l ��]�*��i�u�u�u�w�}��������A9��h_�����b�a�"�0�w�.����	ǹ��T9��\��\��r�r�u�9�2�W�W���Y�Ƽ�9��Q��*���d�
� �d�`��D�ԜY�Ƽ�9��Q��*���d�
� �d�n��D��Y���F���*���3�'�d�
�a�/���Mӑ��]F��R�����'�2�g�`��t�J���^�Ʃ�@�N��U���%�a�7�3�2��C��&���� ^��G]�U���%�a�7�3�2��C�������Q��N�U���u�u�u�2�'�;�(��&����[����*���f�'�2�g�n�u�^��^���V
��d��U���u�%�a�7�1�8�(�������V��N�����7�3�0�
�c�o�(���H����CU�
NךU���u�u�
�
�"�;���&�Г�V��Z�����}�0�
�8��8�(��H���F�G�����_�u�u�u�w��(�������9��h��D��
�f�_�u�w��(�������9��h��D��
�f�i�u�w�}�W���	�ғ�F ��E1�*���'�2�b�a� �8�Wǭ����� 9��P1�L���|�h�r�r�w�1��ԜY���F��1�����
�a�g�
�"�l�Nׁ�J���F��1�����
�a�g�
�"�l�F݁�J���9F�N��U���
�a�u�=�9�u�����ޓ�V��Y�E���u�d�|�0�$�}�W���Y����lR��B����
�a�'�2�`�m�}���Y����Q��R��A��
� �d�d��n�K���Y���F��hZ�� ���'�d�
�a�%�:�@��������h��C���2�g�b�}�~�`�P���Y����l�N��Uʥ�a�7�3�0��i�E݁�����9��d��Uʥ�a�7�3�0��i�Eہ�����9��R�����u�u�u�
��(����Hǹ��l��hY�U���;�}�0�
�:�i����K����O�I�\ʰ�&�u�u�u�w�}��������A9��h\�����a�l�%�n�w�}��������A9��h\�����a�f�%�u�j�W�W���Y�Ƽ�9��Q��*���d�
�0�
�c�}����Q����G��h��*��g�e�u�u�f�t����Y���F���*���3�'�d�
�c�;�(��O����9F���*���3�'�d�
�a�;�(��I����[�N��U���%�a�7�3�2��C��&����R��@��U¦�9�!�%�'�0�o�C���P���A�R��U���u�u�u�%�c�?����&�ғ�9��h_�F���n�u�u�%�c�?����&�ғ�9��h_�B���u�h�_�u�w�}�W���&����V��1�*���
�a�u�=�9�u�����Փ�V��W�E���u�d�|�0�$�}�W���Y����lR��B����
�c�3�
�c�m���Y����lR��B����
�m�3�
�c�i����D���F�N����d�"�0�u�$�1����&����V��^��H��r�u�9�0�]�}�W���Y����Q��R��G���'�2�b�c�]�}�W���&����V��1�*���d�c�
�f�k�}�W���Y����lR��B����
�
�0�
�a�}����Q����G��h��*��l�e�u�u�f�t����Y���F���*���3�'�d�
�o�;�(��M����9F���*���3�'�d�
�g�;�(��A����[�N��U���%�a�7�3�2��E�������P��_��]���
�8�c�'�0�o�@���P���A�R��U���u�u�u�%�c�?����&�ғ�
9��h_�D���n�u�u�%�c�?����&�ғ�9��h_�@���u�h�_�u�w�}�W���&����V��1�����b�c�"�0�w�.����	ǹ��T9��\��\��r�r�u�9�2�W�W���Y�Ƽ�9��Q��*���f�
� �d�a��D�ԜY�Ƽ�9��Q��*���f�
� �d�o��D��Y���F���*���3�'�d�
��8�(��Y����N��[1��؊�0�
�e�g�g�}�W��PӃ��VFǻN��U���
�
� �3�%�l�(�������S��UךU���
�
� �3�%�l�(�������_��N�U���u�u�u�%�c�?����&�ԓ�l��hY�U���;�}�0�
�:�����I���F�_��U���0�_�u�u�w�}�(ہ�����lW��\�� ��m�
�f�_�w�}�(ہ�����lW��Z�� ��l�
�f�i�w�}�W���YӖ��l��Q��D؊�
�0�
�c�w�5��������CU��R	��E��e�u�u�d�~�8����Y���F��hZ�� ���'�d�
�f�1��C���	��ƹF��hZ�� ���'�d�
�`�1��B���	���l�N��Uʥ�a�7�3�0��i����������YN�����8�d�'�2�e�e�_���D����F��D��U���u�u�'�2�o�l�}���Y����Q��R��A��
� �d�d��n�K���Y���F��hZ�� ���'�d�
�
�2��N������@��C��*���
�e�l�e�w�}�F�������9F�N��U���
� �3�'�f��B���&����l��=N��U���
� �3�'�f��@���&����l��S��U���u�u�%�a�5�;����M����V��\�����}�0�
�8�a�/���N����[�I�����u�u�u�u�w�-�C�������R��1��*���e�%�n�u�w�-�C�������R��1��*���a�%�u�h�]�}�W���Y����Q��R��A���'�2�b�g� �8�Wǭ�����9��P1�C���|�h�r�r�w�1��ԜY���F��1�����
�a�f�
�"�l�F؁�J���F��1�����
�a�f�
�"�l�Dށ�J���9F�N��U���
� �3�'�f��(���&����D��F�����%�
�0�
�g�o�G���Y�����RNךU���u�u�
�
�"�;���&�ޓ�F9��Z��F�ߊu�u�
�
�"�;���&����lW��1��U��_�u�u�u�w�/�(���A�ߓ�F��R �����!�%�'�2�e�i�_���D����F��D��U���u�u�%�a�5�;����M�ԓ�V��X�U���%�a�7�3�2��C��&����U��G]��H�ߊu�u�u�u����������@9��P1�Gʢ�0�u�&�9�#�-����K����O�I�\ʰ�&�u�u�u�w�}��������A9��h]�����`�d�%�n�w�}��������A9��hZ�����`�`�%�u�j�W�W���Y�Ƽ�9��Q��*���&�'�2�b�e�*����
����^��E��G��}�|�h�r�p�}����s���F�G1�����0�
�a�a��(�F��&����F�G1�����0�
�a�a�1��D���	���l�N��Uʥ�a�7�3�0��i�E���������YN�����8�f�'�2�e�d�_���D����F��D��U���u�u�%�a�5�;����M�Փ�F9��Z��F�ߊu�u�
�
�"�;���&Ź��lW��1��U��_�u�u�u�w�/�(���A�ߓ�F��R �����!�%�
�0��m�E��Y���O��[�����u�u�u�
��(����Hǹ��A��X����u�
�
� �1�/�Fہ�&���� U��G]��H�ߊu�u�u�u����������9��P1�Gʢ�0�u�&�9�#�-����K����O�I�\ʰ�&�u�u�u�w�}��������A9��hX�� ��g�
�f�_�w�}�(ہ�����lW��1��*��g�%�u�h�]�}�W���Y����Q��R��A���'�2�c�g� �8�Wǭ����� 9��P1�L���|�h�r�r�w�1��ԜY���F��1�����
�a�b�3��n�B���B�����h�����d�
�e�3��h�C���Y���F�N�����3�
�g�
�e�*����
����^��h��*��`�e�u�u�f�t����Y���F���*���3�'�d�
��8�(��B�����h�����d�
�d�3��k�F���Y���F�N�����7�3�0�
�b�d����N����[����*���d�
�0�
�f�h�G���Y�����RNךU���u�u�
�
�"�;���&�֓�F9��Z��F�ߊu�u�
�
�"�;���&�ԓ�F9��V��F��u�u�u�u�w�-�C�������S��h��*��u�=�;�}�2����&����W��^��H��r�u�9�0�]�}�W���Y����Q��R��@��
� �d�e��n�}���Y����Q��R��@��
� �d�d��n�K���Y���F��hZ�� ���'�d�
�
�2��G������@��C��L���2�g�c�}�~�`�P���Y����l�N��Uʥ�a�7�3�0��h�F݁�����9��d��Uʥ�a�7�3�0��h�F؁�����9��R�����u�u�u�0��i�W����έ�l��h�����0�
�8�d��8�(��M����l��^��H��r�u�9�0�]�}�W���Y����Q��R��@��
�0�
�g�l�}�WϮ�M����U��[��M���
�c�l�%�w�`�}���Y���C9��U�����`�d�
�0��o�W����έ�l��h�����0�
�8�d��8�(��L����l��^��H��r�u�9�0�]�}�W���Y����Q��R��@��
� �d�g��n�}���Y����Q��R��@��
� �d�f��n�K���Y���F��hZ�� ���'�d�
�c�%�:�@��������E�����2�&�9�!�'�i����K����C��^�E���u�d�|�0�$�}�W���Y����lR��B����
�m�3�
�a�d���Y����lR��B����
�
� �d�b��D��Y���F�	��*���m�l�%�u�?�3�_���&����
9��P1�C���|�h�r�r�w�1��ԜY���F��1�����
�`�'�2�a�n�}���Y����Q��R��@��
� �d�a��n�K���Y���F��hZ�� ���'�d�
�c�%�:�@��������E�����2�&�9�!�'�n����K����C��^�E���u�d�|�0�$�}�W���Y����lR��B����
�l�3�
�a�k���Y����lR��B����
�d�3�
�a�m����D���F�N��A���3�0�
�`�f�����K�ƻ�V�V�����%�!�
�0��0�Fց�����S��G^�����|�h�r�r�w�1��ԜY���F��1�����
�`�g�
�"�l�C܁�J���F��1�����
�`�g�
�"�l�B؁�J���9F�N��U���
�a�u�=�9�u��������G��R����
�0�
�d�e�-�G���H���F�G�����_�u�u�u�w��(�������9��h��*���n�u�u�%�c�?����&�ӓ� 9��h_�A���u�h�_�u�w�}�W���&����V��1�*���
�`�u�=�9�u��������G��R����
�0�
�d�c�-�G���H���F�G�����_�u�u�u�w��(�������9��h��D���
�f�_�u�w��(�������9��h��D��
�f�i�u�w�}�W���	�ғ�F ��E1�*���'�2�b�f� �8�Wǿ�&����C��P1�����%�`�'�2�e�n�(���&����O�I�\ʰ�&�u�u�u�w�}��������A9��h\�����c�a�%�n�w�}��������A9��h\�����c�m�%�u�j�W�W���Y�Ƽ�9��Q��*���d�
�0�
�b�}����Q����V��G��*���
�8�d�
�2��F���	�֓�GW�N��R��u�9�0�_�w�}�W���&ǹ��U ��h_��Gފ� �d�b�
�d�W�W���&ǹ��U ��h_��G܊� �d�m�
�d�a�W���Y�����h�����d�
�a�'�0�j�Dϩ�����C9��P1�����&�9�!�%�d�/���Hǹ��9��F�U���d�|�0�&�w�}�W���YӖ��l��Q��Dߊ�`�3�
�c�o�-�L���YӖ��l��Q��Dߊ�b�3�
�c�e�-�W��s���F�G1�����0�
�`�d��8�(��Y����N��h��*���!�
�0�
�:�l�(���&����l��h��]���h�r�r�u�;�8�}���Y���C9��U�����`�g�
� �f�e�(��s���C9��U�����`�g�
� �f�d�(��E��ƹF�N�����a�u�=�;��-����	����l��h��DҊ�0�
�d�l�'�m���I���W����ߊu�u�u�u����������@9��P1�L�ߊu�u�
�
�"�;���&�ߓ�F9��X��F��u�u�u�u�w�-�C�������U��h��*��u�=�;�}�'�/����
����V
��Z�*���
�d�g�%�g�4�F��Y���O��[�����u�u�u�
��(����Hƹ��l ��X�*��_�u�u�
��(����Hƹ��l ��Y�*��i�u�u�u�w�}��������A9��h�����b�u�=�;��-����	����l��h��D܊�0�
�d�a�'�m���I���W����ߊu�u�u�u����������_��B1�E܊�f�_�u�u���������� W��B1�Gڊ�f�i�u�u�w�}�WϮ�M����U��]��*���
�b�u�=�9�u��������G��R����
�0�
�d�b�-�G���H���F�G�����_�u�u�u�w��(�������9��h��D��
�f�_�u�w��(�������9��h��D��
�f�i�u�w�}�W���	�ғ�F ��E1�*���0�
�b�u�?�3�_�������C��h��*���d�
�0�
�f�h�������F�_��U���0�_�u�u�w�}�(ہ�����lW��_�� ��g�
�f�_�w�}�(ہ�����lW��]�� ��f�
�f�i�w�}�W���YӖ��l��Q��Dي�
�0�
�b�w�5����	����l��C	�����8�d�
�0��l�C���I����V�
N��R���9�0�_�u�w�}�W���&����V��1�*���d�g�
�f�]�}�W���&����V��1�*���d�a�
�f�k�}�W���Y����lR��B����
�
�0�
�`�}����Q����V��G��*���
�8�d�
�2��F���	�֓�GW�N��R��u�9�0�_�w�}�W���&ǹ��U ��h_��Fي� �d�f�
�d�W�W���&ǹ��U ��h_��Fߊ� �d�a�
�d�a�W���Y�����h�����d�
�
�0��m�W����έ�l��h�����0�
�8�d��8�(��@����l��^��H��r�u�9�0�]�}�W���Y����R��=N��U���
� �3�'�f��A���&����l��S��U���u�u�%�a�5�;����L����V��[�����}�%�'�2�'�.��������Q��R	��D���%�e�<�d�g�}�W��PӃ��VFǻN��U���
�
� �3�%�l�(�������^��UךU���
�
� �3�%�l�(�������T��N�U���u�u�u�%�c�?����&�ӓ�l��hV�U���;�}�%�'�0�-����
����^��h��*��a�%�e�<�f�m�W���H����_��=N��U���u�
�
� �1�/�Fځ�O����Q��h����u�
�
� �1�/�Fځ�A����Q��h�I���u�u�u�u�'�i��������l��R	��E���=�;�}�%�%�:��������l��[�����d�`�%�e�>�l�G���Y�����RNךU���u�u�
�
�"�;���&�ѓ�F9��\��F�ߊu�u�
�
�"�;���&�ߓ�F9�� X��F��u�u�u�u�w�-�C�������S��h��*��u�=�;�}�'�/����
����V
��Z�*���
�d�`�%�g�4�F��Y���O��[�����u�u�u�
��(����Hƹ��l ��Y�*��_�u�u�
��(����Hƹ��U��[�����h�_�u�u�w�}��������l��@��U¦�9�!�%�f�%�:�E��Q���A��N�����u�u�u�u�'�i��������lT��R	��A��u�u�%�a�5�;����L����U�� V�����h�_�u�u�w�}�(ہ�����lW��D1����`�"�0�u�6�����	����@��C��F���2�g�d�
�'�����P���A�R��U���u�u�u�%�c�?����&�ӓ�
9��h_�C���n�u�u�%�c�?����&�ӓ�9��h_�E���u�h�_�u�w�}�W���&����V��1�����m�`�"�0�w�<�(���&����T9��[1�����'�2�g�c��-�(���Q���A��N�����u�u�u�u�'�i��������lR��Q��B���%�n�u�u�'�i��������lR��B1�C܊�f�i�u�u�w�}�WϮ�M����U��[��*���
�a�u�=�9�u��������A��_�]���h�r�r�u�;�8�}���Y���C9��U�����`�f�3�
�b�d���Y����lR��B����
�
� �d�`��D��Y���F�	��*���m�l�%�u�?�3�_���&����9��P1�G���|�h�r�r�w�1��ԜY���F��1�����
�`�`�'�0�k�B�ԜY�Ƽ�9��Q��*���b�3�
�`�g�-�W��s���F�G1�����0�
�`�`�%�:�A��������h��Dي�0�
�d�a�g�}�W��PӃ��VFǻN��U���
�
� �3�%�l�(ف����� 9��d��Uʥ�a�7�3�0��h�O���&����l��S��U���u�u�%�a�5�;����L�ӓ�V�� [�����}�0�
�8�f�����H���F�_��U���0�_�u�u�w�}�(ہ�����lW�� 1��*���e�%�n�_�w�}�ZϮ�N�֓�C9��S1��*���u�&�<�;�'�2����Y��ƹF��hY��*���#�1�<�
�>���������PF��G�����%�b�e�4��1�[Ϯ�N�֓�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(߁�	����O��_�����u�u�u�u�w��(߁�	����l��D��I���
�
�
�%�!�9�}���Y���V
��d��U���u�u�u�%�`�m��������l��R�����e�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��E���
�<�u�&�>�3�������KǻN��*݊�
�;�&�2�6�.���������T��]���
�y�%�b�g�-���	�ѓ�l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`�m�������G��d��U���u�u�u�%�`�m���������h^�U���u�u�0�&�w�}�W���Y�����h^�����2�i�u�
������s���F�R ����_�u�u�;�w�/����B��ƹF�N��B��
�%�#�1�>�����
������T��[���_�u�u�
��m��������l��h�����%�:�u�u�%�>����&Ĺ��l��A��U���
�e�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���4�
�9�|�w�5��ԜY���F�N��B��
�%�#�1�>�����DӖ��lW��V����u�u�u�u�2�.�W���Y���F���*���4�
�9�
�9�.���Y����V��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�N����Z��^	�����;�%�:�0�$�}�Z���YӖ��lW��^ �����&�<�;�%�8�}�W�������C9��^����d�
�'�2�w��(�������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�b�d�
�'�+��������9F�N��U���u�
�
�e�>�����DӖ��lW��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��h�����i�u�
�
�g�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�b�f���������@��V�����'�6�o�%�8�8�Ǯ�N����R��[
����d�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1��Dۊ�%�#�1�|�#�8�W���Y���F���*���4�
�9�
�9�.���Y����W��G1���ߊu�u�u�u�;�8�}���Y���F�G1��Dۊ�%�#�1�<��4�W��	�ѓ�9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&�ד�]9��PN�����u�'�6�&�y�p�}���Y����W��Y1�����&�2�
�'�4�g��������lQ��B��*݊�d�%�0�y�'�j�Fށ�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�d�4��1�^������F�N��U���%�b�d�
�9�.���Y����W��N��U���0�&�u�u�w�}�W���YӖ��lW��^ �����h�%�b�d��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��D؊�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�e�<�(���&����Z��D�����:�u�u�'�4�.�_���&�ԓ�C9��SB��*݊�g�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hY��G���
�9�|�u�?�3�}���Y���F�G1��D؊�%�#�1�<��4�W��	�ѓ�9��h��N���u�u�u�0�$�}�W���Y���F��hY��G���
�9�
�;�$�:�K���&Ĺ��l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����H����l�������%�:�0�&�w�p�W���	�ѓ�9��h��*���<�;�%�:�w�}����
�μ�9��N��B��
�'�2�u���E���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�b�d�
�%�!�9�^Ϫ���ƹF�N��U���
�
�g�<��4�W��	�ѓ�]ǻN��U���9�0�_�u�w�}�W���Y����T��Y1����u�
�
�g�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��F���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�b�d��-��������T9��D��*���6�o�%�:�2�.����H����l��N��B��
�%�#�1�'�8�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F�� 1�*���#�1�|�!�2�}�W���Y���F��hY��F���
�9�
�;�$�:�K���&Ĺ��l��A�����u�u�u�9�2�W�W���Y���F�� 1�*���#�1�<�
�>�}�JϮ�N����R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(؁�J����@��V�����'�6�&�{�z�W�W���&Ĺ��l��D�����2�
�'�6�m�-����
ۖ��lW����*���%�0�y�%�`�l�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�f�4�
�;�t�W������F�N��Uʥ�b�d�
�;�$�:�K���&Ĺ��l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ� 9��h��U��%�b�d�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F�� 1�*���#�1�<�
�>�}����Ӗ��P��N����u�
�
�a�6���������l��^	�����u�u�'�6�$�u�(؁�M����E
����*���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h_�����9�|�u�=�9�W�W���Y���F�� 1�*���#�1�<�
�>�}�JϮ�N����R��[
�U���u�u�0�&�w�}�W���Y�����h_�����9�
�;�&�0�a�W���&�ғ�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@��&����Z��D��ʥ�:�0�&�u�z�}�WϮ�N����Z��^	�����;�%�:�u�w�/����Q����R�G1��Dފ�'�2�u�
��i������ƹF��R	�����u�u�u�3��<�(���
����T��N�����d�
�%�#�3�t����Y���F�N��U���
�a�<�
�>�}�JϮ�N����9F�N��U���0�_�u�u�w�}�W���&Ĺ��l��D��I���
�
�a�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h_�����9�
�;�&�0�<����Y����V��C�U���%�b�d�
�'�+����&����R��P �����o�%�:�0�$�-�@��&����_�G1��Dߊ�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��[�����1�|�!�0�w�}�W���Y�����h_�����9�
�;�&�0�a�W���&�ӓ�C9��SUךU���u�u�9�0�]�}�W���Y���C9��[�����1�<�
�<�w�`����Hƹ��l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������TF��D��U���6�&�{�x�]�}�W���&�ӓ�]9��P1�����
�'�6�o�'�2����	�ѓ�J��hY��@���0�y�%�b�f��������F��P��U���u�u�<�u��-��������Z��S��*݊�`�4�
�9�~�}����s���F�N�����d�
�;�&�0�a�W���&����F�N�����u�u�u�u�w�}�WϮ�N����Z��^	��Hʥ�b�d�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��1��*���
�;�&�2�6�.��������@H�d��Uʥ�b�d�4�
�;���������Z��G��U���'�6�&�}���(������C9��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ѓ�l��A��\ʡ�0�u�u�u�w�}�W���	�ѓ�l��A�����<�u�h�%�`�l������ƹF�N�����_�u�u�u�w�}�W���&¹��l��h�����i�u�
�
��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�
�;�$�:�����Ƽ�\��D@��X���u�%�b�d�>�����
����l��TN����0�&�%�b�f�}�(؁�&����F�� 1�����9�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&¹��l��G�����_�u�u�u�w�}�W���&¹��l��R�����d�_�u�u�w�}����s���F�N�����d�<�
�<�w�`����H����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�
�'�+����&����R��P �����&�{�x�_�w�}�(؁�&����_��Y1�����&�2�
�'�4�g��������lQ��h�����u�
�
�
�'�+������ƹF��R	�����u�u�u�3��<�(���
����T��N�����g�4�
�9�~�}����s���F�N�����g�4�
�9��3����E�Ƽ�9��V����u�u�u�u�2�.�W���Y���F���*؊�%�#�1�<��4�W��	�ѓ�l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����K����@��V�����'�6�&�{�z�W�W���&Ĺ��Z��^	�����;�%�:�u�w�/����Q����J��hY��*���2�u�
�
��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*؊�%�#�1�|�#�8�W���Y���F���*؊�;�&�2�i�w��(��Y���F��[�����u�u�u�u�w��(݁�����Z�G1��G���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�N�Փ�C9��S1��*���u�&�<�;�'�2����Y��ƹF��hY��*���#�1�<�
�>���������PF��G�����%�b�f�4��1�[Ϯ�N�Փ�C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(܁�	����O��_�����u�u�u�u�w��(܁�	����l��D��I���
�
�
�%�!�9�}���Y���V
��d��U���u�u�u�%�`�n��������l��R�����f�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��F���
�<�u�&�>�3�������KǻN��*݊�
�;�&�2�6�.���������T��]���
�y�%�b�d�-���	�ѓ�l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�`�n�������G��d��U���u�u�u�%�`�n���������h]�U���u�u�0�&�w�}�W���Y�����h]�����2�i�u�
������s���F�R ����_�u�u�;�w�/����B��ƹF�N��B���4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�b�c�<�(���&����Z��D�����:�u�u�'�4�.�_���&ǹ��l��N��B���4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������hZ�����1�|�!�0�w�}�W���Y�����hZ�����1�<�
�<�w�`����M����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��V�����;�&�2�i�w��(ہ�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
������Ӈ��Z��G�����u�x�u�u�'�j�C���&����R��P �����o�%�:�0�$�-�@��Y����9��R	����a�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��V�����u�=�;�_�w�}�W���Y�Ƽ�9��^ �����h�%�b�a�]�}�W���Y����l�N��U���u�%�b�a�>�����DӖ��lR��E�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u���(�������]9��PN�����u�'�6�&�y�p�}���Y����9��h��*���&�2�4�&�0�����CӖ��P����*ߊ�%�#�1�u���(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�b�`�6�����Y����l�N��U���u�%�b�`�6���������Z�G1��@���
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�%�!�9���������h[�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lS��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��1��*���
�&�<�;�'�2�W�������@N�� 1�U���
�
�'�2�w��(ځ�	����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�;�$�:�K���&Ĺ��9F�N��U���0�_�u�u�w�}�W���&Ĺ��Z��^	��Hʥ�b�`�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lQ��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�`�k��������lQ��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&Ĺ��R��[
��U���;�_�u�u�w�}�W���&Ĺ��R��[
�����2�i�u�
���������F�N�����u�u�u�u�w�}����O����E
��^ �����h�%�b�c�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�b�c�<�
�>�}����Ӗ��P��N����u�
�
�
�9�.����
����C��T�����&�}�
�
�{�-�@���	������hX�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����O����E
��N�����u�u�u�u�w�}����O����@��S��*݊�n�u�u�u�w�8����Y���F�N��*݊�
�;�&�2�k�}�(؁�&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�b�b�4��1�(���
����@��YN�����&�u�x�u�w�-�@�������W9��h��*���<�;�%�:�w�}����
�μ�9��V�����%�b�b�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*݊�
�%�#�1�~�)����Y���F�N��*݊�
�%�#�1�>�����DӖ��lQ��G1���ߊu�u�u�u�;�8�}���Y���F�G1��B���
�9�
�;�$�:�K���&Ĺ��R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(؁�&����Z��D��ʥ�:�0�&�u�z�}�WϮ�N�ѓ�]9��P1�����
�'�6�o�'�2����	�ѓ�F�� 1�����y�%�b�b�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��B���
�9�|�u�?�3�}���Y���F�G1��B���
�<�u�h�'�j�@�ԜY���F��D��U���u�u�u�u�'�j�@���&����[��hY��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&˹��l��h�����4�&�2�u�%�>���T���F�� 1�����9�
�;�&�0�<����&����\��E�����
�
�
�%�!�9�W���&˹��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�j�O���&����F��R ��U���u�u�u�u�'�j�O���&����Z��^	��Hʥ�b�m�4�
�;�f�W���Y����_��=N��U���u�u�u�
����������@��S��*݊�
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hY��*���&�2�4�&�0�}����
���l�N��B���<�
�<�
�$�4��������C��R�����m�u�
�
��/����&Ĺ��R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
����������[��=N��U���u�u�u�
���������C9��UךU���u�u�9�0�]�}�W���Y���C9��1��*���u�h�%�b�o�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*ӊ�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��-��������T9��D��*���6�o�%�:�2�.����@����E
����*ӊ�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��1��*���|�u�=�;�]�}�W���Y���C9��1��*���
�;�&�2�k�}�(؁�&����_��N��U���0�&�u�u�w�}�W���YӖ��l_��G1�����
�<�u�h�'�j�N���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�b�n�4�(���Y����T��E�����x�_�u�u���(���
����@��Y1�����u�'�6�&���(��	�ѓ�l��PB��*݊�
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l_��G1�����!�0�u�u�w�}�W���YӖ��l_��Y1����u�
�
�n�w�}�W�������9F�N��U���u�
�
�
�9�.���Y����
9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n�m��������l�������%�:�0�&�w�p�W���	�ߓ�l��A�����<�
�&�<�9�-����Y����V��G1��E���
�9�y�%�n�m��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�'�+��������9F�N��U���u�
�
�
�'�+����&����[��hW��*���#�1�_�u�w�}�W������F�N��Uʥ�l�e�4�
�;��������C9��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��h��U���<�;�%�:�2�.�W��Y����l_��h�����4�&�2�
�%�>�MϮ�������h^����e�%�0�y�'�d�G���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�l�e�4�
�;�t�W������F�N��Uʥ�l�e�<�
�>�}�JϮ�@����F�N�����u�u�u�u�w�}�WϮ�@�֓�]9��PN�U���
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�e�4�
�;���������Z��G��U���'�6�&�}���G���&������h_�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lW��V�����u�=�;�_�w�}�W���Y�Ƽ�
9��h�����<�
�<�u�j�-�N��&����_��N��U���0�&�u�u�w�}�W���YӖ��lW��V�����;�&�2�i�w��(�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n�l�(���
����@��YN�����&�u�x�u�w�-�N��&����Z��D�����:�u�u�'�4�.�_���&���C9��^�����u�
�
�e�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��Dڊ�%�#�1�|�#�8�W���Y���F���*���<�
�<�u�j�-�N��B���F����ߊu�u�u�u�w�}�(ց�I����@��S��*ӊ�e�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��lW��V�����;�&�2�4�$�:�W�������K��N�����d�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�n�l�(������C9��_�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����W��G1�����!�0�u�u�w�}�W���YӖ��lW��V�����;�&�2�i�w��(�������W]ǻN��U���9�0�_�u�w�}�W���Y����W��G1�����
�<�u�h�'�d�Fށ�	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��l�����ƭ�@�������{�x�_�u�w��(�������T9��D��*���6�o�%�:�2�.����H����l_��1�����%�l�d�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hW��D���
�9�|�u�?�3�}���Y���F�G1��Dۊ�;�&�2�i�w��(��s���F�R��U���u�u�u�u�w�-�N��&����Z�
N��L��
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����T��G1�����
�<�u�&�>�3�������KǻN��*ӊ�g�4�
�9��3��������]9��X��U���6�&�}�
��o��������l_��1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ߓ�9��h��\���=�;�_�u�w�}�W���Y����T��G1�����
�<�u�h�'�d�F݁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ߓ�9��h��*���&�2�i�u���E���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�l�f�����Ӈ��Z��G�����u�x�u�u�'�d�F݁�����l��^	�����u�u�'�6�$�u�(ց�K�Ƽ�
9��h�����
�
�g�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�*���#�1�|�!�2�}�W���Y���F��hW��G���
�<�u�h�'�d�F��Y���F��[�����u�u�u�u�w��(�������TF���*���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ߓ� 9��h��*���&�2�4�&�0�}����
���l�N��L��
�%�#�1�>�����
����l��TN����0�&�%�l�f������Ƽ�
9��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ʹ��l��A��\ʡ�0�u�u�u�w�}�W���	�ߓ� 9��h��*���&�2�i�u���D���&����9F�N��U���0�_�u�u�w�}�W���&ʹ��l��A�����<�u�h�%�n�l�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�d�4�(���Y����T��E�����x�_�u�u���D���&����R��P �����o�%�:�0�$�-�N��UӖ��lW��G��Yʥ�l�d�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h_�����9�|�u�=�9�W�W���Y���F��1�*���&�2�i�u���D�ԜY���F��D��U���u�u�u�u�'�d�F܁�����Z�G1��Dي�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ʹ��l��A�����<�u�&�<�9�-����
���9F���*���4�
�9�
�9�.����
����C��T�����&�}�
�
�c�<�(���UӖ��lW��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�@����R��[
��U���;�_�u�u�w�}�W���&ʹ��l��A�����<�u�h�%�n�l�(�������F�N�����u�u�u�u�w�}�WϮ�@����R��[
�����2�i�u�
��i��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�l�d��3��������]F��X�����x�u�u�%�n�l�(���
����@��Y1�����u�'�6�&���(��Y����R��E��U���
�a�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��Z�����1�|�!�0�w�}�W���Y�����h_�����<�u�h�%�n�l�L���Y�����RNךU���u�u�u�u���C���&����[��hW��A���0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�@����R��[
�����2�4�&�2�w�/����W���F�G1��Dߊ�%�#�1�<��4�(�������A	��N�����&�%�l�d��-����Y����S��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&�ӓ�C9��SG�����u�u�u�u�w�}�WϮ�@����R��[
�����2�i�u�
��h������ƹF�N�����_�u�u�u�w�}�W���&�ӓ�C9��S1��*���u�h�%�l�f���������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�
�`�>�����
������T��[���_�u�u�
��h��������@��h����%�:�0�&�'�d�F��	�ߓ�9��R	����d�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����l_��1��*���|�u�=�;�]�}�W���Y���C9��[�����2�i�u�
��h�}���Y���V
��d��U���u�u�u�%�n�l�(���
���F��1�*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&¹��l��h�����4�&�2�u�%�>���T���F��1�����9�
�;�&�0�<����&����\��E�����
�
�
�%�!�9�W���&¹��l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�d�F���&����F��R ��U���u�u�u�u�'�d�F���&����Z��^	��Hʥ�l�d�4�
�;�f�W���Y����_��=N��U���u�u�u�
����������@��S��*ӊ�
�%�#�1�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��hW��*���&�2�4�&�0�}����
���l�N��L���<�
�<�
�$�4��������C��R�����d�u�
�
��/����&ʹ��R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
����������[��=N��U���u�u�u�
���������C9��UךU���u�u�9�0�]�}�W���Y���C9��1��*���u�h�%�l�f�-���Y���F��Y
�����u�u�0�1�'�2����s���F���*؊�%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��-��������T9��D��*���6�o�%�:�2�.����K����E
����*؊�%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��1��*���|�u�=�;�]�}�W���Y���C9��1��*���
�;�&�2�k�}�(ց�&����_��N��U���0�&�u�u�w�}�W���YӖ��lT��G1�����
�<�u�h�'�d�E���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�l�e�4�(���Y����T��E�����x�_�u�u���(���
����@��Y1�����u�'�6�&���(��	�ߓ�l��PB��*ӊ�
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��lT��G1�����!�0�u�u�w�}�W���YӖ��lT��Y1����u�
�
�n�w�}�W�������9F�N��U���u�
�
�
�9�.���Y����9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�n�n��������l�������%�:�0�&�w�p�W���	�ߓ�l��A�����<�
�&�<�9�-����Y����V��G1��F���
�9�y�%�n�n��������V�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�
�'�+��������9F�N��U���u�
�
�
�'�+����&����[��hW��*���#�1�_�u�w�}�W������F�N��Uʥ�l�f�4�
�;��������C9��1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y���� 9��h��U���<�;�%�:�2�.�W��Y����l_��h�����4�&�2�
�%�>�MϮ�������h]����f�%�0�y�'�d�D���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�l�f�4�
�;�t�W������F�N��Uʥ�l�f�<�
�>�}�JϮ�@����F�N�����u�u�u�u�w�}�WϮ�@�Փ�]9��PN�U���
�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�
9��V�����;�&�2�4�$�:�W�������K��N�����a�4�
�9��3��������]9��X��U���6�&�}�
�������Ƽ�
9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�@�ғ�C9��SG�����u�u�u�u�w�}�WϮ�@�ғ�C9��S1��*���u�h�%�l�c�<�(���B���F����ߊu�u�u�u�w�}�(ց�&����_��Y1����u�
�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�
�;�&�0�<����Y����V��C�U���%�l�a�<��4�(�������A	��N�����&�%�l�a�w��(ہ����C9��1��*���|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}�(ց�&����_����ߊu�u�u�u�w�}�(ց�&����Z�
N��L��_�u�u�u�w�1��ԜY���F�N��L���<�
�<�u�j�-�N���	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�
�%�!�9�����ƭ�@�������{�x�_�u�w��(ځ�	����l��D�����2�
�'�6�m�-����
ۖ��lS��G1�����
�
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��L���4�
�9�|�w�5��ԜY���F�N��L���4�
�9�
�9�.���Y����9��h��N���u�u�u�0�$�}�W���Y���F��hW��*���#�1�<�
�>�}�JϮ�@�ӓ�C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�N�������TF��D��U���6�&�{�x�]�}�W���&ƹ��l��h�����%�:�u�u�%�>����&ʹ����h[�����u�
�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��hW��*���#�1�|�!�2�}�W���Y���F��hW��*���&�2�i�u���L���Y�����RNךU���u�u�u�u���(���
���F��1�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p����O����E
��^ �����&�<�;�%�8�8����T�����hX�����1�<�
�<��.����	����	F��X��¥�l�c�4�
�;�q����O����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u���(��������YNךU���u�u�u�u���(�������]9��PN�U���
�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�l�a�<�(���&����Z�
N��L���4�
�9�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1�����<�u�&�<�9�-����
���9F���*܊�;�&�2�4�$�:�(�������A	��D��*ӊ�y�%�l�c�'�8�[Ϯ�@�Г�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�l�a�<�(���P�Ƹ�V�N��U���u�u�%�l�a�4�(���Y����l_��d��U���u�0�&�u�w�}�W���Y����l_��h�����i�u�
�
��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1��B���
�9�
�;�$�:�����Ƽ�\��D@��X���u�%�l�b�6���������l��^	�����u�u�'�6�$�u�(ց�&����_�G1��B���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����l_��h�����|�!�0�u�w�}�W���Y����l_��h�����<�
�<�u�j�-�N�������W]ǻN��U���9�0�_�u�w�}�W���Y����9��h��*���&�2�i�u���(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
��3��������]F��X�����x�u�u�%�n�j��������@��h����%�:�0�&�'�d�@���&ʹ��C��N��L���4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����9��h��\���=�;�_�u�w�}�W���Y����9��h��U��%�l�b�_�w�}�W������F�N��U���%�l�b�<��4�W��	�ߓ�l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
����������@��V�����'�6�&�{�z�W�W���&ʹ��R��[
�����2�4�&�2��/���	����@��hW��*���#�1�u�
����������TOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�l�m�4��1�^������F�N��U���%�l�m�4��1�(���
���F��1�����9�n�u�u�w�}����Y���F�N��U���
�
�%�#�3�4�(���Y����l_��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ߓ�l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�
9��^ �����&�<�;�%�8�}�W�������C9��B��*ӊ�
�'�2�u���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�%�#�3�t����Y���F�N��U���
�
�;�&�0�a�W���&��ƹF�N�����_�u�u�u�w�}�W���&˹��l��R�����m�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l_��G1�����
�<�u�&�>�3�������KǻN��*ӊ�
�%�#�1�>�����
����l��TN����0�&�%�l�n�<�(���UӖ��l_��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&ʹ��l��G�����_�u�u�u�w�}�W���&ʹ��l��h�����i�u�
�
��-����s���F�R��U���u�u�u�u�w�-�N�������W9��h��U��%�l�l�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����l�<�
�<�w�.����	����@�CךU���
�
�
�;�$�:��������\������}�
�
�y�'�d�N�������l_��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�N�������WO�C��U���u�u�u�u�w�-�N�������TF���*��u�u�u�u�2�.�W���Y���F���*ӊ�;�&�2�i�w��(ց�����F�N�����<�n�_�u�w�3�W�������9l�N�����%�e�3�
�g�j����D���F�N��L���<�
�<�u�?�3�_���&����l ��Y�����|�h�r�r�w�1��ԜY���F��[1��ӊ� �d�f�
�d�W�W�������CW��Q��E���%�u�h�_�w�}�W���&ʹ��l��D�����u�&�9�!�'����@����O�I�\ʰ�&�u�u�u�w�}��������l ��^�*��_�u�u�0��0�F݁�����9��R�����u�u�u�
��o�����ƻ�V�D�����
� �m�`�'�u�^��^���V
��d��U���u�&�9�!�'�l����I�ғ� ]ǻN�����8�d�
� �f�j�(��E���F��R �����<��'��8��(ށ�Kù��U��Y�����u�%�6�;�#�1�C��Y����D��d��Uʦ�9�!�%�a�1��G���	���D��������9�
�:��2����H����l��B1�Bۊ�g�h�4�
�8�.�(���&����_��^�����u�0�
�8�f����Aʹ��Z�_�����u�<�
�<��/�;���&ƹ��T��C1��*��d�%�u�u�'�>�����ғ�F��D��E��u�u�&�9�#�-�A���&����l��S��D���=�;�}��;���������lW��^��*���d�b�
�g�j�<�(���
����9�������w�_�u�u�2����&����V��G\��H���w�"�0�u�>���������C9��1�E���3�
�e�d�'�}�W�������l
��h,�����u�e�n�u�w�.����	�ޓ�F9��Y��G��u�d�u�=�9�u�;���&����	��h[��*��
�
� �d�`��E������]��[��1���9�0�w�w�]�}�W���&����
9��h_�F���u�h�w�w� �8�WǷ�&����\��X��@���e�e�!�3��m�F���Y�ƭ�l��D��ފ�|�0�&�u�g�f�W���
����^��Q��Mߊ�g�i�u�d�w�5��������l^��h�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����8�g�
� �f�n�(��E��ƹF�N��*ӊ�
�;�&�2� �8�Wǭ�����U��B1�B݊�g�e�u�u�f�t����Y���F���*���<�
�<�n�w�}��������l ��\�*��i�u�u�u�w�}����L����@��@��U¦�9�!�%�a�1��G���	����[�I�����u�u�u�u�w�.����	�֓�F9��W��F�ߊu�u�0�
�:�o�(���H����CU�
NךU���u�u�
�
��3����������h��Dߊ� �d�m�
�e�m�W���H����_��=N��U���u�0�
�8�e����Mƹ��l�N�����%�f�3�
�e�d����D���F�N��L���<�
�<�u�?�3�_���&����9��h_�@���}�|�h�r�p�}����s���F�D�����g�3�
�g�e�-�L���Yӕ��l��Z�� ��c�
�f�i�w�}�W���YӖ��lW��^ �����=�;�}�0��0�F؁�����9��^��H��r�u�9�0�]�}�W���Y����G��1��*��l�%�n�u�w�.����	�ӓ�F9�� ]��F��u�u�u�u�w�-�N��&����Z��_��]���
�8�d�
�"�l�G؁�K���F�G�����_�u�u�u�w�8�(���Kǹ��lW��1��N���u�&�9�!�'����H����[�L�����}�8�
� �o�l����Y����\��h��*���0�&�u�e�l�}�Wϭ����� 9��hV�*��i�u�d�u�?�3�_���&����W��N�����:�&�
�#��t����Y���9F���*���a�3�
�c��o�K���H�ƻ�V�C�����`�
�d�h�6�����&����O��[��W���_�u�u�0��0�B���&����l��S��U���u�u�%�l�e�4�(���Y����N��[1�����
�`�
�g�g�}�W��PӃ��VFǻN��U���
�
�a�<��4�L���Yӕ��l��1��*��
�g�i�u�f�}����Q����U��_��D��4�
�:�&��+�(�������V�=N��U���
�8�b�3��m�D���Y���F�N�����a�<�
�<�w�5��������CT��B1�D���}�|�h�r�p�}����s���F�D�����
� �d�d��n�}���Y����G��h��M���%�u�h�w�u�*��������F9��1��U���%�6�;�!�;�i�6������D��N�����!�%�
� �f�n�(��E��ƹF�N��*ӊ�
�;�&�2� �8�Wǭ�����9��hV�*��e�u�u�d�~�8����Y���F��R�����3�
�e�f�'�f�W���
����^��B1�@���u�h�w�w� �8�WǪ�	����S��G_��U���6�;�!�9�c�o�W�������l�N�����
�`�
�d�k�}�;���&����	��h[����� �m�g�%��}�W�������V�=��U���4�n�