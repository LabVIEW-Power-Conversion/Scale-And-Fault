-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��E���M����l��X��Fئ�f�
�u�&�w�}�������9F�N��U���u�u�u�u�m�4�������]ǻN��U��� �
���w�g�������F��=N��U���u�<�e����MϷ�����\�\�U���u�u�1� ���#���Y����T��S��G���u�|�_�u�w�2����Y���F��[��U���;�u�!�
�8�4�L���Y�����R��U���u�!�
�:�>�f�W���Y����VF�T�����!�
�:�<�l�}�W���Yӂ��F���U���
�:�<�
�2�)�Ǻ�ù��w2��N�����u�|�_�u�w�}�W�������\��D�����6�#�6�:��2����=�����Y��E�ߊu�u�n�0�3�8����B���P��R�����'�=�:�u��o�E����֓�Z��G1���
�u�&�u�w�p�Z��T���K�C�X���:�%�;�;�w�p�Z��T���K�C�X���u�6�8�:�2�)���H����U9��V�����%�e�;�
�$��EϷ�s���F�G��U�ߊu�u�u�u�w�}�(���
����E��SN��U���u�;�u�!��2���Y���F�N��*���&�4�!�4�6�}�W���Cӏ����h�����0�!�'�f�w�2����I��ƹF�N��U���
�-�&�'�$�1�(������	����*���<�n�u�u�w�}�W�������@9��D��*���!�u�o�:�#�.��������V��EF�U���;�:�e�_�w�}�W���B����������;�n�u�u�z�p�Z��T���K�C�U���4�u�<�;�;�p�Z��T���K�C�U���&�2�4�u��+����Y�ƿ�W9��P�����u�<�;�9�6�)����Y����G��X	��*���!�'�f�u�8�3���B�����Y�����4�<�u�o�$�9�������F��P ��U���1�!�u�u�w�)�(�������P��]����!�u�|�_�w�}����ӂ��9��Q_��U���
�:�<�
�2�)�Ǻ�ù��w2��N�����u�|�_�0�>�W�W���T���K�C�X���x�x��&�6�)�������K�C�X���x�_�u�u��o�E����֓�C9��C��*ڊ�:�1�%�f��}�W���	����GF��\�1ޔ�
�
�%�&�#�;�(߁�����lU��N�����u�4�u�_�w�}�W���&����l��A�����u�u�k�4�#�<���Y���F��h�����!�4�4�u�w�}�J���&����RJǻN��U���
�-�&�'�$�1�(������F��C�����u�u�u�u�:�<��������l��C��H���
�1�!�_�w�}�L�ԜY���K�C�X���x�x�x�x��.�������K�C�X���x�x�x�_�w�}�(������F�UךU���
�1�!�u�k�}����&����{K��S�����u�k�r�r�w�5��������Q��S��U���e����f�9� ���Y���A��G�����1�;�
� �f�`�_Ϻ�ù��w2��N�����u�u�k�r�p�t�W���ӂ��9��Q_�U���1� �u�u�w�`��������9F�C�X���x�x�x�x�z�p�Z�������Q��R��X���x�x�x�x�z�p�Z���YӖ��P��F�����0�<�_�u�w�}�W�������E����U���u�u�d�u�?�3�W���Y���F��QN��U���d�u�=�;�w�}�W���Y���F��^ �����u�h�1�;�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R����1�4�6�<�2�)���