-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�<����V��1�����c�g�'�8�>�}�W�������Z�N��U���u�u�8�8�#�-�W���Cӕ��Z��S�����>�n�_�u�w�}�W���Y����G�N��U���0�0�u�h�d�f�}���Y���F�V�����u�u�u�;�2�8�W��M��ƹF�N��U���0�
�<�0�w�}�W�������	[�d��U���u�u�u�%�%�}�}���Y���F��S�U���o�<�u�!��2����������S��Dʱ�"�!�u�|�w�}�W���Y����VV�N��U���;�&�1�9�0�>�W���Y���F��N��U���u�u� �u�#�����&����\��@����1�"�!�u�~�W�W���Y���R��N��U��<�u�!�
�8�4�(�������D��_C����!�u�|�u�w�}�W���YӅ��F�N��U���&�1�9�2�4�}�W���Y�����N��U���u�;�&�1�;�:��������W��C��U���;�:�e�n�]�}�W���Y�ƻ�F�N��Oʼ�u�!�
�:�>�f�}���Y���F��N��U���o�:�!�&�3�1��������AN��^
��X���:�;�:�e�l�}�W���Y����_�N��U��<�u�!�
�8�4�W���Y����9�������u�_�4�6�>�8����Y����\ ��+�B��3�e�4�,�g�k�E���ӏ��9l��P ��U���'�
�8�u�w�)�(�������P�������d�1�"�!�w�t�W������R��1����&�1�9�2�4�+����Q����G�
�����e�n�_�,�2�0��������@F��E��]���:�8�8�&�-�p�^ϱ�Y����_	��T1�����u�1�<�!�z�}�������l��V��U���<�7�0�'�:�g��������l��C�����u�,�
�4�$�$���
����T]�V�����0�&�;�'�:�)����Ӕ��\��V�����<�u�7�:�<�/�������Q����*���9�u�u�!�>�:�}�������VF��Z1�����:�u�4�u�w�<����ӏ��^��C��N��!�<� �0���!���7����t/��r<��0����u�u�!�>�:�}�����9l��Z��*���0�&�2�4�3�m�W���������E^�����<�_�u�u�w�9�߁������E^�XǦ�;�=�&�&�#�<��������9F�N��������������I���^��D��X���!�0�_�u�w�}�W�������l��R��]���0�&�h�u�g�t�}���Y�Ʃ�@�N��U���u�u�1�'��0�W������l�N�����<�n�x�&�9�5��������_��h�����%�:�0�&�]�-��������P��h^����0�&�}�9�~�}�������F��F��Ͱ�0�!�4�1�4�6�J���^�Ƹ�VǻN��U���3�}�0�u�w�l�^Ϫ���ƹF�N��U���e�i�u�4���!���-������E^�����n�_�u�u�w�}�������F��SN��N��1�%�:�0�$�W��������P��h	�����o�%�:�0�$�u����P���T��N��Uʴ�1�d�!�%�k�}����B����J��R��U���;�9�!�
�1�W�W���Y���p)��h'��0���}�1�'�|�i�0����������Yd��U���u�u�u�1�%�����D�Σ�[��S�R��n�u�u�u�2�.�W���Y���F�V
��D���%�i�u�1�%�f�W���YӃ����=C�����0�<�u�'�9�1����������T��N���
�0�:�,�6�>����CӖ��P��F�����_�0�<�u�w�}��������E����U���u�u�d�|�#�8�}���Y���Z �T�H��r�u�=�;�]�}�W���Y���Z �@�H��r�u�=�;�]�}�W���Y���F�E��6���
�����9�ށ����	[��U��U���u�u�u�u�2�9���Y���F�N��D��u�4�}����#���+ۇ��AW��Z��N�ߊu�u�u�u�9�}��ԜY�Ʃ�WF��d��ʥ�:�0�&�_�]�3�W���B����Z��E��0���_�&�u���.��������P��V����!�!�u�`�f�j�F߸�I����lV��\�����u�2�;�'�4�u�W���Y����R��^
��U������u�j�n�L���Y���'��E��'���0�o�����M���O���F�N�����&�<�!�u�w��2���Y���]ǻN�����}�u�u�u�w�/����Cӯ��`2��{!��6�ߊu�u�u�u�;�}�W���*����|!��d��U���u�4�1�0�$�}�W���*����|!��h8��!����1�0�&�>�)�W���Y����g)�UךU���u�u�0�u�w��$���5����l�N��Uʤ�u�u� �u���8���&����|4��V�����u�u�u����G��Y���F��S
����o��u����>���<����'��E��"���=�x�d�� �	�W���s���F�T�Oʜ�u��
���f�W���Y����VW�'��&������_�w�}�W���H����}F��s1��2������}�6�<����Y����w)��c!��\�ߊu�u�u�u�f�g�8���*����|!��h8��!����!��1�?�p�FϚ�.����O�=��U���<�,�_�4�4�4�����ƭ�P��QN��0���e�
�
�%��(��Y��ƹF��X�����u�`�d�b�f�;�G��� �֓�T��V�����u�u�u�%�%�}�}���Y���F�T��Oʜ�u��
���f�W���Y���F��S
��U���������!���6��ƹF�N��U���0�u�u����;���:���F�N��Uʤ�u�u� �u���8���&����|4��N��U���u�u�4�1�f�g�>���-����t/��a+��:��u�u�u�u�w�}���Cӯ��`2��{!��6�ߊu�u�u�u�w�}�F��0�Ɵ�w9��p'��#����n�u�u�w�}�W������/��d:��9����_�u�u�w�}�W���H����f2��c*��:���
����l�}�Wϻ�Ӆ��C	��Y����0�<�_�u�w�h�F���HÀ��l��h^��E؊�4�
�u�u�4�0����Ӌ��_��^��E���,�e�c�g�%�0�W���	����^��d��U���u�6�>�h�w�1�[���Y�����E^��Kʴ�1�0�&�y�w�}�W������F��BךU���u�u�e�h�w�m�}���Y���R��N��U���'�&�d�_�w�}�W��������d��U���u�1�u�k�3�q�W���Y����VW�	N��D�ߊu�u�u�u�f�`�W��B���WF��T�����'�n�_�